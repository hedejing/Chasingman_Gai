module bkg_tile_table(
	addr,
	q
);
input  [12: 0] addr;
output reg [ 2: 0] q;

always @(*)
	case(addr)
	13'd0: q = 3'b000;
	13'd1: q = 3'b000;
	13'd2: q = 3'b000;
	13'd3: q = 3'b000;
	13'd4: q = 3'b000;
	13'd5: q = 3'b000;
	13'd6: q = 3'b000;
	13'd7: q = 3'b000;
	13'd8: q = 3'b000;
	13'd9: q = 3'b000;
	13'd10: q = 3'b000;
	13'd11: q = 3'b000;
	13'd12: q = 3'b000;
	13'd13: q = 3'b000;
	13'd14: q = 3'b000;
	13'd15: q = 3'b000;
	13'd16: q = 3'b000;
	13'd17: q = 3'b000;
	13'd18: q = 3'b000;
	13'd19: q = 3'b000;
	13'd20: q = 3'b000;
	13'd21: q = 3'b000;
	13'd22: q = 3'b000;
	13'd23: q = 3'b000;
	13'd24: q = 3'b000;
	13'd25: q = 3'b000;
	13'd26: q = 3'b000;
	13'd27: q = 3'b000;
	13'd28: q = 3'b000;
	13'd29: q = 3'b000;
	13'd30: q = 3'b000;
	13'd31: q = 3'b000;
	13'd32: q = 3'b000;
	13'd33: q = 3'b000;
	13'd34: q = 3'b000;
	13'd35: q = 3'b000;
	13'd36: q = 3'b000;
	13'd37: q = 3'b000;
	13'd38: q = 3'b000;
	13'd39: q = 3'b000;
	13'd40: q = 3'b000;
	13'd41: q = 3'b000;
	13'd42: q = 3'b000;
	13'd43: q = 3'b000;
	13'd44: q = 3'b000;
	13'd45: q = 3'b000;
	13'd46: q = 3'b000;
	13'd47: q = 3'b000;
	13'd48: q = 3'b000;
	13'd49: q = 3'b000;
	13'd50: q = 3'b000;
	13'd51: q = 3'b000;
	13'd52: q = 3'b000;
	13'd53: q = 3'b000;
	13'd54: q = 3'b000;
	13'd55: q = 3'b000;
	13'd56: q = 3'b000;
	13'd57: q = 3'b000;
	13'd58: q = 3'b000;
	13'd59: q = 3'b000;
	13'd60: q = 3'b000;
	13'd61: q = 3'b000;
	13'd62: q = 3'b000;
	13'd63: q = 3'b000;
	13'd64: q = 3'b000;
	13'd65: q = 3'b000;
	13'd66: q = 3'b000;
	13'd67: q = 3'b000;
	13'd68: q = 3'b000;
	13'd69: q = 3'b000;
	13'd70: q = 3'b000;
	13'd71: q = 3'b000;
	13'd72: q = 3'b000;
	13'd73: q = 3'b000;
	13'd74: q = 3'b000;
	13'd75: q = 3'b000;
	13'd76: q = 3'b000;
	13'd77: q = 3'b000;
	13'd78: q = 3'b000;
	13'd79: q = 3'b000;
	13'd80: q = 3'b000;
	13'd81: q = 3'b000;
	13'd82: q = 3'b000;
	13'd83: q = 3'b000;
	13'd84: q = 3'b000;
	13'd85: q = 3'b000;
	13'd86: q = 3'b000;
	13'd87: q = 3'b000;
	13'd88: q = 3'b000;
	13'd89: q = 3'b000;
	13'd90: q = 3'b000;
	13'd91: q = 3'b000;
	13'd92: q = 3'b000;
	13'd93: q = 3'b000;
	13'd94: q = 3'b000;
	13'd95: q = 3'b000;
	13'd96: q = 3'b000;
	13'd97: q = 3'b000;
	13'd98: q = 3'b000;
	13'd99: q = 3'b000;
	13'd100: q = 3'b000;
	13'd101: q = 3'b000;
	13'd102: q = 3'b000;
	13'd103: q = 3'b000;
	13'd104: q = 3'b000;
	13'd105: q = 3'b000;
	13'd106: q = 3'b000;
	13'd107: q = 3'b000;
	13'd108: q = 3'b000;
	13'd109: q = 3'b000;
	13'd110: q = 3'b000;
	13'd111: q = 3'b000;
	13'd112: q = 3'b000;
	13'd113: q = 3'b000;
	13'd114: q = 3'b000;
	13'd115: q = 3'b000;
	13'd116: q = 3'b000;
	13'd117: q = 3'b000;
	13'd118: q = 3'b000;
	13'd119: q = 3'b000;
	13'd120: q = 3'b000;
	13'd121: q = 3'b000;
	13'd122: q = 3'b000;
	13'd123: q = 3'b000;
	13'd124: q = 3'b000;
	13'd125: q = 3'b000;
	13'd126: q = 3'b000;
	13'd127: q = 3'b000;
	13'd128: q = 3'b000;
	13'd129: q = 3'b000;
	13'd130: q = 3'b000;
	13'd131: q = 3'b000;
	13'd132: q = 3'b000;
	13'd133: q = 3'b000;
	13'd134: q = 3'b000;
	13'd135: q = 3'b000;
	13'd136: q = 3'b000;
	13'd137: q = 3'b000;
	13'd138: q = 3'b000;
	13'd139: q = 3'b000;
	13'd140: q = 3'b000;
	13'd141: q = 3'b000;
	13'd142: q = 3'b000;
	13'd143: q = 3'b000;
	13'd144: q = 3'b000;
	13'd145: q = 3'b000;
	13'd146: q = 3'b000;
	13'd147: q = 3'b000;
	13'd148: q = 3'b000;
	13'd149: q = 3'b000;
	13'd150: q = 3'b000;
	13'd151: q = 3'b000;
	13'd152: q = 3'b000;
	13'd153: q = 3'b000;
	13'd154: q = 3'b000;
	13'd155: q = 3'b000;
	13'd156: q = 3'b000;
	13'd157: q = 3'b000;
	13'd158: q = 3'b000;
	13'd159: q = 3'b000;
	13'd160: q = 3'b000;
	13'd161: q = 3'b000;
	13'd162: q = 3'b000;
	13'd163: q = 3'b000;
	13'd164: q = 3'b000;
	13'd165: q = 3'b000;
	13'd166: q = 3'b000;
	13'd167: q = 3'b000;
	13'd168: q = 3'b000;
	13'd169: q = 3'b000;
	13'd170: q = 3'b000;
	13'd171: q = 3'b000;
	13'd172: q = 3'b000;
	13'd173: q = 3'b000;
	13'd174: q = 3'b000;
	13'd175: q = 3'b000;
	13'd176: q = 3'b000;
	13'd177: q = 3'b000;
	13'd178: q = 3'b000;
	13'd179: q = 3'b000;
	13'd180: q = 3'b000;
	13'd181: q = 3'b000;
	13'd182: q = 3'b000;
	13'd183: q = 3'b000;
	13'd184: q = 3'b000;
	13'd185: q = 3'b000;
	13'd186: q = 3'b000;
	13'd187: q = 3'b000;
	13'd188: q = 3'b000;
	13'd189: q = 3'b000;
	13'd190: q = 3'b000;
	13'd191: q = 3'b000;
	13'd192: q = 3'b000;
	13'd193: q = 3'b000;
	13'd194: q = 3'b000;
	13'd195: q = 3'b000;
	13'd196: q = 3'b000;
	13'd197: q = 3'b000;
	13'd198: q = 3'b000;
	13'd199: q = 3'b000;
	13'd200: q = 3'b000;
	13'd201: q = 3'b000;
	13'd202: q = 3'b000;
	13'd203: q = 3'b000;
	13'd204: q = 3'b000;
	13'd205: q = 3'b000;
	13'd206: q = 3'b000;
	13'd207: q = 3'b000;
	13'd208: q = 3'b000;
	13'd209: q = 3'b000;
	13'd210: q = 3'b000;
	13'd211: q = 3'b000;
	13'd212: q = 3'b000;
	13'd213: q = 3'b000;
	13'd214: q = 3'b000;
	13'd215: q = 3'b000;
	13'd216: q = 3'b000;
	13'd217: q = 3'b000;
	13'd218: q = 3'b000;
	13'd219: q = 3'b000;
	13'd220: q = 3'b000;
	13'd221: q = 3'b000;
	13'd222: q = 3'b000;
	13'd223: q = 3'b000;
	13'd224: q = 3'b000;
	13'd225: q = 3'b000;
	13'd226: q = 3'b000;
	13'd227: q = 3'b000;
	13'd228: q = 3'b000;
	13'd229: q = 3'b000;
	13'd230: q = 3'b000;
	13'd231: q = 3'b000;
	13'd232: q = 3'b000;
	13'd233: q = 3'b000;
	13'd234: q = 3'b000;
	13'd235: q = 3'b000;
	13'd236: q = 3'b000;
	13'd237: q = 3'b000;
	13'd238: q = 3'b000;
	13'd239: q = 3'b000;
	13'd240: q = 3'b000;
	13'd241: q = 3'b000;
	13'd242: q = 3'b000;
	13'd243: q = 3'b000;
	13'd244: q = 3'b000;
	13'd245: q = 3'b000;
	13'd246: q = 3'b000;
	13'd247: q = 3'b000;
	13'd248: q = 3'b000;
	13'd249: q = 3'b000;
	13'd250: q = 3'b000;
	13'd251: q = 3'b000;
	13'd252: q = 3'b000;
	13'd253: q = 3'b000;
	13'd254: q = 3'b000;
	13'd255: q = 3'b000;
	13'd256: q = 3'b000;
	13'd257: q = 3'b000;
	13'd258: q = 3'b000;
	13'd259: q = 3'b000;
	13'd260: q = 3'b000;
	13'd261: q = 3'b000;
	13'd262: q = 3'b000;
	13'd263: q = 3'b000;
	13'd264: q = 3'b000;
	13'd265: q = 3'b000;
	13'd266: q = 3'b000;
	13'd267: q = 3'b000;
	13'd268: q = 3'b000;
	13'd269: q = 3'b000;
	13'd270: q = 3'b000;
	13'd271: q = 3'b000;
	13'd272: q = 3'b000;
	13'd273: q = 3'b000;
	13'd274: q = 3'b000;
	13'd275: q = 3'b000;
	13'd276: q = 3'b000;
	13'd277: q = 3'b000;
	13'd278: q = 3'b000;
	13'd279: q = 3'b000;
	13'd280: q = 3'b000;
	13'd281: q = 3'b000;
	13'd282: q = 3'b000;
	13'd283: q = 3'b000;
	13'd284: q = 3'b000;
	13'd285: q = 3'b000;
	13'd286: q = 3'b000;
	13'd287: q = 3'b000;
	13'd288: q = 3'b000;
	13'd289: q = 3'b000;
	13'd290: q = 3'b000;
	13'd291: q = 3'b000;
	13'd292: q = 3'b000;
	13'd293: q = 3'b000;
	13'd294: q = 3'b000;
	13'd295: q = 3'b000;
	13'd296: q = 3'b000;
	13'd297: q = 3'b000;
	13'd298: q = 3'b000;
	13'd299: q = 3'b000;
	13'd300: q = 3'b000;
	13'd301: q = 3'b000;
	13'd302: q = 3'b000;
	13'd303: q = 3'b000;
	13'd304: q = 3'b000;
	13'd305: q = 3'b000;
	13'd306: q = 3'b000;
	13'd307: q = 3'b000;
	13'd308: q = 3'b000;
	13'd309: q = 3'b000;
	13'd310: q = 3'b000;
	13'd311: q = 3'b000;
	13'd312: q = 3'b000;
	13'd313: q = 3'b000;
	13'd314: q = 3'b000;
	13'd315: q = 3'b000;
	13'd316: q = 3'b000;
	13'd317: q = 3'b000;
	13'd318: q = 3'b000;
	13'd319: q = 3'b000;
	13'd320: q = 3'b000;
	13'd321: q = 3'b000;
	13'd322: q = 3'b000;
	13'd323: q = 3'b000;
	13'd324: q = 3'b000;
	13'd325: q = 3'b000;
	13'd326: q = 3'b000;
	13'd327: q = 3'b000;
	13'd328: q = 3'b000;
	13'd329: q = 3'b000;
	13'd330: q = 3'b000;
	13'd331: q = 3'b000;
	13'd332: q = 3'b000;
	13'd333: q = 3'b000;
	13'd334: q = 3'b000;
	13'd335: q = 3'b000;
	13'd336: q = 3'b000;
	13'd337: q = 3'b000;
	13'd338: q = 3'b000;
	13'd339: q = 3'b000;
	13'd340: q = 3'b000;
	13'd341: q = 3'b000;
	13'd342: q = 3'b000;
	13'd343: q = 3'b000;
	13'd344: q = 3'b000;
	13'd345: q = 3'b000;
	13'd346: q = 3'b000;
	13'd347: q = 3'b000;
	13'd348: q = 3'b000;
	13'd349: q = 3'b000;
	13'd350: q = 3'b000;
	13'd351: q = 3'b000;
	13'd352: q = 3'b000;
	13'd353: q = 3'b000;
	13'd354: q = 3'b000;
	13'd355: q = 3'b000;
	13'd356: q = 3'b000;
	13'd357: q = 3'b000;
	13'd358: q = 3'b000;
	13'd359: q = 3'b000;
	13'd360: q = 3'b000;
	13'd361: q = 3'b000;
	13'd362: q = 3'b000;
	13'd363: q = 3'b000;
	13'd364: q = 3'b000;
	13'd365: q = 3'b000;
	13'd366: q = 3'b000;
	13'd367: q = 3'b000;
	13'd368: q = 3'b000;
	13'd369: q = 3'b000;
	13'd370: q = 3'b000;
	13'd371: q = 3'b000;
	13'd372: q = 3'b000;
	13'd373: q = 3'b000;
	13'd374: q = 3'b000;
	13'd375: q = 3'b000;
	13'd376: q = 3'b000;
	13'd377: q = 3'b000;
	13'd378: q = 3'b000;
	13'd379: q = 3'b000;
	13'd380: q = 3'b000;
	13'd381: q = 3'b000;
	13'd382: q = 3'b000;
	13'd383: q = 3'b000;
	13'd384: q = 3'b000;
	13'd385: q = 3'b000;
	13'd386: q = 3'b000;
	13'd387: q = 3'b000;
	13'd388: q = 3'b000;
	13'd389: q = 3'b000;
	13'd390: q = 3'b000;
	13'd391: q = 3'b000;
	13'd392: q = 3'b000;
	13'd393: q = 3'b000;
	13'd394: q = 3'b000;
	13'd395: q = 3'b000;
	13'd396: q = 3'b000;
	13'd397: q = 3'b000;
	13'd398: q = 3'b000;
	13'd399: q = 3'b000;
	13'd400: q = 3'b000;
	13'd401: q = 3'b000;
	13'd402: q = 3'b000;
	13'd403: q = 3'b000;
	13'd404: q = 3'b000;
	13'd405: q = 3'b000;
	13'd406: q = 3'b000;
	13'd407: q = 3'b000;
	13'd408: q = 3'b000;
	13'd409: q = 3'b000;
	13'd410: q = 3'b000;
	13'd411: q = 3'b000;
	13'd412: q = 3'b000;
	13'd413: q = 3'b000;
	13'd414: q = 3'b000;
	13'd415: q = 3'b000;
	13'd416: q = 3'b000;
	13'd417: q = 3'b000;
	13'd418: q = 3'b000;
	13'd419: q = 3'b000;
	13'd420: q = 3'b000;
	13'd421: q = 3'b000;
	13'd422: q = 3'b000;
	13'd423: q = 3'b000;
	13'd424: q = 3'b000;
	13'd425: q = 3'b000;
	13'd426: q = 3'b000;
	13'd427: q = 3'b000;
	13'd428: q = 3'b000;
	13'd429: q = 3'b000;
	13'd430: q = 3'b000;
	13'd431: q = 3'b000;
	13'd432: q = 3'b000;
	13'd433: q = 3'b000;
	13'd434: q = 3'b000;
	13'd435: q = 3'b000;
	13'd436: q = 3'b000;
	13'd437: q = 3'b000;
	13'd438: q = 3'b000;
	13'd439: q = 3'b000;
	13'd440: q = 3'b000;
	13'd441: q = 3'b000;
	13'd442: q = 3'b000;
	13'd443: q = 3'b000;
	13'd444: q = 3'b000;
	13'd445: q = 3'b000;
	13'd446: q = 3'b000;
	13'd447: q = 3'b000;
	13'd448: q = 3'b000;
	13'd449: q = 3'b000;
	13'd450: q = 3'b000;
	13'd451: q = 3'b000;
	13'd452: q = 3'b000;
	13'd453: q = 3'b000;
	13'd454: q = 3'b000;
	13'd455: q = 3'b000;
	13'd456: q = 3'b000;
	13'd457: q = 3'b000;
	13'd458: q = 3'b000;
	13'd459: q = 3'b000;
	13'd460: q = 3'b000;
	13'd461: q = 3'b000;
	13'd462: q = 3'b000;
	13'd463: q = 3'b000;
	13'd464: q = 3'b000;
	13'd465: q = 3'b000;
	13'd466: q = 3'b000;
	13'd467: q = 3'b000;
	13'd468: q = 3'b000;
	13'd469: q = 3'b000;
	13'd470: q = 3'b000;
	13'd471: q = 3'b000;
	13'd472: q = 3'b000;
	13'd473: q = 3'b000;
	13'd474: q = 3'b000;
	13'd475: q = 3'b000;
	13'd476: q = 3'b000;
	13'd477: q = 3'b000;
	13'd478: q = 3'b000;
	13'd479: q = 3'b000;
	13'd480: q = 3'b000;
	13'd481: q = 3'b000;
	13'd482: q = 3'b000;
	13'd483: q = 3'b000;
	13'd484: q = 3'b000;
	13'd485: q = 3'b000;
	13'd486: q = 3'b000;
	13'd487: q = 3'b000;
	13'd488: q = 3'b000;
	13'd489: q = 3'b000;
	13'd490: q = 3'b000;
	13'd491: q = 3'b000;
	13'd492: q = 3'b000;
	13'd493: q = 3'b000;
	13'd494: q = 3'b000;
	13'd495: q = 3'b000;
	13'd496: q = 3'b000;
	13'd497: q = 3'b000;
	13'd498: q = 3'b000;
	13'd499: q = 3'b000;
	13'd500: q = 3'b000;
	13'd501: q = 3'b000;
	13'd502: q = 3'b000;
	13'd503: q = 3'b000;
	13'd504: q = 3'b000;
	13'd505: q = 3'b000;
	13'd506: q = 3'b000;
	13'd507: q = 3'b000;
	13'd508: q = 3'b000;
	13'd509: q = 3'b000;
	13'd510: q = 3'b000;
	13'd511: q = 3'b000;
	13'd512: q = 3'b000;
	13'd513: q = 3'b000;
	13'd514: q = 3'b000;
	13'd515: q = 3'b000;
	13'd516: q = 3'b000;
	13'd517: q = 3'b000;
	13'd518: q = 3'b000;
	13'd519: q = 3'b000;
	13'd520: q = 3'b000;
	13'd521: q = 3'b000;
	13'd522: q = 3'b000;
	13'd523: q = 3'b000;
	13'd524: q = 3'b000;
	13'd525: q = 3'b000;
	13'd526: q = 3'b000;
	13'd527: q = 3'b000;
	13'd528: q = 3'b000;
	13'd529: q = 3'b000;
	13'd530: q = 3'b000;
	13'd531: q = 3'b000;
	13'd532: q = 3'b000;
	13'd533: q = 3'b000;
	13'd534: q = 3'b000;
	13'd535: q = 3'b000;
	13'd536: q = 3'b000;
	13'd537: q = 3'b000;
	13'd538: q = 3'b000;
	13'd539: q = 3'b000;
	13'd540: q = 3'b000;
	13'd541: q = 3'b000;
	13'd542: q = 3'b000;
	13'd543: q = 3'b000;
	13'd544: q = 3'b000;
	13'd545: q = 3'b000;
	13'd546: q = 3'b000;
	13'd547: q = 3'b000;
	13'd548: q = 3'b000;
	13'd549: q = 3'b000;
	13'd550: q = 3'b000;
	13'd551: q = 3'b000;
	13'd552: q = 3'b000;
	13'd553: q = 3'b000;
	13'd554: q = 3'b000;
	13'd555: q = 3'b000;
	13'd556: q = 3'b000;
	13'd557: q = 3'b000;
	13'd558: q = 3'b000;
	13'd559: q = 3'b000;
	13'd560: q = 3'b000;
	13'd561: q = 3'b000;
	13'd562: q = 3'b000;
	13'd563: q = 3'b000;
	13'd564: q = 3'b000;
	13'd565: q = 3'b000;
	13'd566: q = 3'b000;
	13'd567: q = 3'b000;
	13'd568: q = 3'b000;
	13'd569: q = 3'b000;
	13'd570: q = 3'b000;
	13'd571: q = 3'b000;
	13'd572: q = 3'b000;
	13'd573: q = 3'b000;
	13'd574: q = 3'b000;
	13'd575: q = 3'b000;
	13'd576: q = 3'b000;
	13'd577: q = 3'b000;
	13'd578: q = 3'b000;
	13'd579: q = 3'b000;
	13'd580: q = 3'b000;
	13'd581: q = 3'b000;
	13'd582: q = 3'b000;
	13'd583: q = 3'b000;
	13'd584: q = 3'b000;
	13'd585: q = 3'b000;
	13'd586: q = 3'b000;
	13'd587: q = 3'b000;
	13'd588: q = 3'b000;
	13'd589: q = 3'b000;
	13'd590: q = 3'b000;
	13'd591: q = 3'b000;
	13'd592: q = 3'b000;
	13'd593: q = 3'b000;
	13'd594: q = 3'b000;
	13'd595: q = 3'b000;
	13'd596: q = 3'b000;
	13'd597: q = 3'b000;
	13'd598: q = 3'b000;
	13'd599: q = 3'b000;
	13'd600: q = 3'b000;
	13'd601: q = 3'b000;
	13'd602: q = 3'b000;
	13'd603: q = 3'b000;
	13'd604: q = 3'b000;
	13'd605: q = 3'b000;
	13'd606: q = 3'b000;
	13'd607: q = 3'b000;
	13'd608: q = 3'b000;
	13'd609: q = 3'b000;
	13'd610: q = 3'b000;
	13'd611: q = 3'b000;
	13'd612: q = 3'b000;
	13'd613: q = 3'b000;
	13'd614: q = 3'b000;
	13'd615: q = 3'b000;
	13'd616: q = 3'b000;
	13'd617: q = 3'b000;
	13'd618: q = 3'b000;
	13'd619: q = 3'b000;
	13'd620: q = 3'b000;
	13'd621: q = 3'b000;
	13'd622: q = 3'b000;
	13'd623: q = 3'b000;
	13'd624: q = 3'b000;
	13'd625: q = 3'b000;
	13'd626: q = 3'b000;
	13'd627: q = 3'b000;
	13'd628: q = 3'b000;
	13'd629: q = 3'b000;
	13'd630: q = 3'b000;
	13'd631: q = 3'b000;
	13'd632: q = 3'b000;
	13'd633: q = 3'b000;
	13'd634: q = 3'b000;
	13'd635: q = 3'b000;
	13'd636: q = 3'b000;
	13'd637: q = 3'b000;
	13'd638: q = 3'b000;
	13'd639: q = 3'b000;
	13'd640: q = 3'b000;
	13'd641: q = 3'b000;
	13'd642: q = 3'b000;
	13'd643: q = 3'b000;
	13'd644: q = 3'b000;
	13'd645: q = 3'b000;
	13'd646: q = 3'b000;
	13'd647: q = 3'b000;
	13'd648: q = 3'b000;
	13'd649: q = 3'b000;
	13'd650: q = 3'b000;
	13'd651: q = 3'b000;
	13'd652: q = 3'b000;
	13'd653: q = 3'b000;
	13'd654: q = 3'b000;
	13'd655: q = 3'b000;
	13'd656: q = 3'b000;
	13'd657: q = 3'b000;
	13'd658: q = 3'b000;
	13'd659: q = 3'b000;
	13'd660: q = 3'b000;
	13'd661: q = 3'b000;
	13'd662: q = 3'b000;
	13'd663: q = 3'b000;
	13'd664: q = 3'b000;
	13'd665: q = 3'b000;
	13'd666: q = 3'b000;
	13'd667: q = 3'b000;
	13'd668: q = 3'b000;
	13'd669: q = 3'b000;
	13'd670: q = 3'b000;
	13'd671: q = 3'b000;
	13'd672: q = 3'b000;
	13'd673: q = 3'b000;
	13'd674: q = 3'b000;
	13'd675: q = 3'b000;
	13'd676: q = 3'b000;
	13'd677: q = 3'b000;
	13'd678: q = 3'b000;
	13'd679: q = 3'b000;
	13'd680: q = 3'b000;
	13'd681: q = 3'b000;
	13'd682: q = 3'b000;
	13'd683: q = 3'b000;
	13'd684: q = 3'b000;
	13'd685: q = 3'b000;
	13'd686: q = 3'b000;
	13'd687: q = 3'b000;
	13'd688: q = 3'b000;
	13'd689: q = 3'b000;
	13'd690: q = 3'b000;
	13'd691: q = 3'b000;
	13'd692: q = 3'b000;
	13'd693: q = 3'b000;
	13'd694: q = 3'b000;
	13'd695: q = 3'b000;
	13'd696: q = 3'b000;
	13'd697: q = 3'b000;
	13'd698: q = 3'b000;
	13'd699: q = 3'b000;
	13'd700: q = 3'b000;
	13'd701: q = 3'b000;
	13'd702: q = 3'b000;
	13'd703: q = 3'b000;
	13'd704: q = 3'b000;
	13'd705: q = 3'b000;
	13'd706: q = 3'b000;
	13'd707: q = 3'b000;
	13'd708: q = 3'b000;
	13'd709: q = 3'b000;
	13'd710: q = 3'b000;
	13'd711: q = 3'b000;
	13'd712: q = 3'b000;
	13'd713: q = 3'b000;
	13'd714: q = 3'b000;
	13'd715: q = 3'b000;
	13'd716: q = 3'b000;
	13'd717: q = 3'b000;
	13'd718: q = 3'b000;
	13'd719: q = 3'b000;
	13'd720: q = 3'b000;
	13'd721: q = 3'b000;
	13'd722: q = 3'b000;
	13'd723: q = 3'b000;
	13'd724: q = 3'b000;
	13'd725: q = 3'b000;
	13'd726: q = 3'b000;
	13'd727: q = 3'b000;
	13'd728: q = 3'b000;
	13'd729: q = 3'b000;
	13'd730: q = 3'b000;
	13'd731: q = 3'b000;
	13'd732: q = 3'b000;
	13'd733: q = 3'b000;
	13'd734: q = 3'b000;
	13'd735: q = 3'b000;
	13'd736: q = 3'b000;
	13'd737: q = 3'b000;
	13'd738: q = 3'b000;
	13'd739: q = 3'b000;
	13'd740: q = 3'b000;
	13'd741: q = 3'b000;
	13'd742: q = 3'b000;
	13'd743: q = 3'b000;
	13'd744: q = 3'b000;
	13'd745: q = 3'b000;
	13'd746: q = 3'b000;
	13'd747: q = 3'b000;
	13'd748: q = 3'b000;
	13'd749: q = 3'b000;
	13'd750: q = 3'b000;
	13'd751: q = 3'b000;
	13'd752: q = 3'b000;
	13'd753: q = 3'b000;
	13'd754: q = 3'b000;
	13'd755: q = 3'b000;
	13'd756: q = 3'b000;
	13'd757: q = 3'b000;
	13'd758: q = 3'b000;
	13'd759: q = 3'b000;
	13'd760: q = 3'b000;
	13'd761: q = 3'b000;
	13'd762: q = 3'b000;
	13'd763: q = 3'b000;
	13'd764: q = 3'b000;
	13'd765: q = 3'b000;
	13'd766: q = 3'b000;
	13'd767: q = 3'b000;
	13'd768: q = 3'b000;
	13'd769: q = 3'b000;
	13'd770: q = 3'b000;
	13'd771: q = 3'b000;
	13'd772: q = 3'b000;
	13'd773: q = 3'b000;
	13'd774: q = 3'b000;
	13'd775: q = 3'b000;
	13'd776: q = 3'b000;
	13'd777: q = 3'b000;
	13'd778: q = 3'b000;
	13'd779: q = 3'b000;
	13'd780: q = 3'b000;
	13'd781: q = 3'b000;
	13'd782: q = 3'b000;
	13'd783: q = 3'b000;
	13'd784: q = 3'b000;
	13'd785: q = 3'b000;
	13'd786: q = 3'b000;
	13'd787: q = 3'b000;
	13'd788: q = 3'b000;
	13'd789: q = 3'b000;
	13'd790: q = 3'b000;
	13'd791: q = 3'b000;
	13'd792: q = 3'b000;
	13'd793: q = 3'b000;
	13'd794: q = 3'b000;
	13'd795: q = 3'b000;
	13'd796: q = 3'b000;
	13'd797: q = 3'b000;
	13'd798: q = 3'b000;
	13'd799: q = 3'b000;
	13'd800: q = 3'b000;
	13'd801: q = 3'b000;
	13'd802: q = 3'b000;
	13'd803: q = 3'b000;
	13'd804: q = 3'b000;
	13'd805: q = 3'b000;
	13'd806: q = 3'b000;
	13'd807: q = 3'b000;
	13'd808: q = 3'b000;
	13'd809: q = 3'b000;
	13'd810: q = 3'b000;
	13'd811: q = 3'b000;
	13'd812: q = 3'b000;
	13'd813: q = 3'b000;
	13'd814: q = 3'b000;
	13'd815: q = 3'b000;
	13'd816: q = 3'b000;
	13'd817: q = 3'b000;
	13'd818: q = 3'b000;
	13'd819: q = 3'b000;
	13'd820: q = 3'b000;
	13'd821: q = 3'b000;
	13'd822: q = 3'b000;
	13'd823: q = 3'b000;
	13'd824: q = 3'b000;
	13'd825: q = 3'b000;
	13'd826: q = 3'b000;
	13'd827: q = 3'b000;
	13'd828: q = 3'b000;
	13'd829: q = 3'b000;
	13'd830: q = 3'b000;
	13'd831: q = 3'b000;
	13'd832: q = 3'b000;
	13'd833: q = 3'b000;
	13'd834: q = 3'b000;
	13'd835: q = 3'b000;
	13'd836: q = 3'b000;
	13'd837: q = 3'b000;
	13'd838: q = 3'b000;
	13'd839: q = 3'b000;
	13'd840: q = 3'b000;
	13'd841: q = 3'b000;
	13'd842: q = 3'b000;
	13'd843: q = 3'b000;
	13'd844: q = 3'b000;
	13'd845: q = 3'b000;
	13'd846: q = 3'b000;
	13'd847: q = 3'b000;
	13'd848: q = 3'b000;
	13'd849: q = 3'b000;
	13'd850: q = 3'b000;
	13'd851: q = 3'b000;
	13'd852: q = 3'b000;
	13'd853: q = 3'b000;
	13'd854: q = 3'b000;
	13'd855: q = 3'b000;
	13'd856: q = 3'b000;
	13'd857: q = 3'b000;
	13'd858: q = 3'b000;
	13'd859: q = 3'b000;
	13'd860: q = 3'b000;
	13'd861: q = 3'b000;
	13'd862: q = 3'b000;
	13'd863: q = 3'b000;
	13'd864: q = 3'b000;
	13'd865: q = 3'b000;
	13'd866: q = 3'b000;
	13'd867: q = 3'b000;
	13'd868: q = 3'b000;
	13'd869: q = 3'b000;
	13'd870: q = 3'b000;
	13'd871: q = 3'b000;
	13'd872: q = 3'b000;
	13'd873: q = 3'b000;
	13'd874: q = 3'b000;
	13'd875: q = 3'b000;
	13'd876: q = 3'b000;
	13'd877: q = 3'b000;
	13'd878: q = 3'b000;
	13'd879: q = 3'b000;
	13'd880: q = 3'b000;
	13'd881: q = 3'b000;
	13'd882: q = 3'b000;
	13'd883: q = 3'b000;
	13'd884: q = 3'b000;
	13'd885: q = 3'b000;
	13'd886: q = 3'b000;
	13'd887: q = 3'b000;
	13'd888: q = 3'b000;
	13'd889: q = 3'b000;
	13'd890: q = 3'b000;
	13'd891: q = 3'b000;
	13'd892: q = 3'b000;
	13'd893: q = 3'b000;
	13'd894: q = 3'b000;
	13'd895: q = 3'b000;
	13'd896: q = 3'b000;
	13'd897: q = 3'b000;
	13'd898: q = 3'b000;
	13'd899: q = 3'b000;
	13'd900: q = 3'b000;
	13'd901: q = 3'b000;
	13'd902: q = 3'b000;
	13'd903: q = 3'b000;
	13'd904: q = 3'b000;
	13'd905: q = 3'b000;
	13'd906: q = 3'b000;
	13'd907: q = 3'b000;
	13'd908: q = 3'b000;
	13'd909: q = 3'b000;
	13'd910: q = 3'b000;
	13'd911: q = 3'b000;
	13'd912: q = 3'b000;
	13'd913: q = 3'b000;
	13'd914: q = 3'b000;
	13'd915: q = 3'b000;
	13'd916: q = 3'b000;
	13'd917: q = 3'b000;
	13'd918: q = 3'b000;
	13'd919: q = 3'b000;
	13'd920: q = 3'b000;
	13'd921: q = 3'b000;
	13'd922: q = 3'b000;
	13'd923: q = 3'b000;
	13'd924: q = 3'b000;
	13'd925: q = 3'b000;
	13'd926: q = 3'b000;
	13'd927: q = 3'b000;
	13'd928: q = 3'b000;
	13'd929: q = 3'b000;
	13'd930: q = 3'b000;
	13'd931: q = 3'b000;
	13'd932: q = 3'b000;
	13'd933: q = 3'b000;
	13'd934: q = 3'b000;
	13'd935: q = 3'b000;
	13'd936: q = 3'b000;
	13'd937: q = 3'b000;
	13'd938: q = 3'b000;
	13'd939: q = 3'b000;
	13'd940: q = 3'b000;
	13'd941: q = 3'b000;
	13'd942: q = 3'b000;
	13'd943: q = 3'b000;
	13'd944: q = 3'b000;
	13'd945: q = 3'b000;
	13'd946: q = 3'b000;
	13'd947: q = 3'b000;
	13'd948: q = 3'b000;
	13'd949: q = 3'b000;
	13'd950: q = 3'b000;
	13'd951: q = 3'b000;
	13'd952: q = 3'b000;
	13'd953: q = 3'b000;
	13'd954: q = 3'b000;
	13'd955: q = 3'b000;
	13'd956: q = 3'b000;
	13'd957: q = 3'b000;
	13'd958: q = 3'b000;
	13'd959: q = 3'b000;
	13'd960: q = 3'b000;
	13'd961: q = 3'b000;
	13'd962: q = 3'b000;
	13'd963: q = 3'b000;
	13'd964: q = 3'b000;
	13'd965: q = 3'b000;
	13'd966: q = 3'b000;
	13'd967: q = 3'b000;
	13'd968: q = 3'b000;
	13'd969: q = 3'b000;
	13'd970: q = 3'b000;
	13'd971: q = 3'b000;
	13'd972: q = 3'b000;
	13'd973: q = 3'b000;
	13'd974: q = 3'b000;
	13'd975: q = 3'b000;
	13'd976: q = 3'b000;
	13'd977: q = 3'b000;
	13'd978: q = 3'b000;
	13'd979: q = 3'b000;
	13'd980: q = 3'b000;
	13'd981: q = 3'b000;
	13'd982: q = 3'b000;
	13'd983: q = 3'b000;
	13'd984: q = 3'b000;
	13'd985: q = 3'b000;
	13'd986: q = 3'b000;
	13'd987: q = 3'b000;
	13'd988: q = 3'b000;
	13'd989: q = 3'b000;
	13'd990: q = 3'b000;
	13'd991: q = 3'b000;
	13'd992: q = 3'b000;
	13'd993: q = 3'b000;
	13'd994: q = 3'b000;
	13'd995: q = 3'b000;
	13'd996: q = 3'b000;
	13'd997: q = 3'b000;
	13'd998: q = 3'b000;
	13'd999: q = 3'b000;
	13'd1000: q = 3'b000;
	13'd1001: q = 3'b000;
	13'd1002: q = 3'b000;
	13'd1003: q = 3'b000;
	13'd1004: q = 3'b000;
	13'd1005: q = 3'b000;
	13'd1006: q = 3'b000;
	13'd1007: q = 3'b000;
	13'd1008: q = 3'b000;
	13'd1009: q = 3'b000;
	13'd1010: q = 3'b000;
	13'd1011: q = 3'b000;
	13'd1012: q = 3'b000;
	13'd1013: q = 3'b000;
	13'd1014: q = 3'b000;
	13'd1015: q = 3'b000;
	13'd1016: q = 3'b000;
	13'd1017: q = 3'b000;
	13'd1018: q = 3'b000;
	13'd1019: q = 3'b000;
	13'd1020: q = 3'b000;
	13'd1021: q = 3'b000;
	13'd1022: q = 3'b000;
	13'd1023: q = 3'b000;
	13'd1024: q = 3'b011;
	13'd1025: q = 3'b011;
	13'd1026: q = 3'b111;
	13'd1027: q = 3'b111;
	13'd1028: q = 3'b111;
	13'd1029: q = 3'b111;
	13'd1030: q = 3'b111;
	13'd1031: q = 3'b111;
	13'd1032: q = 3'b111;
	13'd1033: q = 3'b111;
	13'd1034: q = 3'b111;
	13'd1035: q = 3'b111;
	13'd1036: q = 3'b111;
	13'd1037: q = 3'b111;
	13'd1038: q = 3'b111;
	13'd1039: q = 3'b111;
	13'd1040: q = 3'b111;
	13'd1041: q = 3'b111;
	13'd1042: q = 3'b111;
	13'd1043: q = 3'b111;
	13'd1044: q = 3'b111;
	13'd1045: q = 3'b111;
	13'd1046: q = 3'b111;
	13'd1047: q = 3'b111;
	13'd1048: q = 3'b111;
	13'd1049: q = 3'b111;
	13'd1050: q = 3'b111;
	13'd1051: q = 3'b111;
	13'd1052: q = 3'b111;
	13'd1053: q = 3'b111;
	13'd1054: q = 3'b000;
	13'd1055: q = 3'b000;
	13'd1056: q = 3'b011;
	13'd1057: q = 3'b011;
	13'd1058: q = 3'b111;
	13'd1059: q = 3'b111;
	13'd1060: q = 3'b111;
	13'd1061: q = 3'b111;
	13'd1062: q = 3'b111;
	13'd1063: q = 3'b111;
	13'd1064: q = 3'b111;
	13'd1065: q = 3'b111;
	13'd1066: q = 3'b111;
	13'd1067: q = 3'b111;
	13'd1068: q = 3'b111;
	13'd1069: q = 3'b111;
	13'd1070: q = 3'b111;
	13'd1071: q = 3'b111;
	13'd1072: q = 3'b111;
	13'd1073: q = 3'b111;
	13'd1074: q = 3'b111;
	13'd1075: q = 3'b111;
	13'd1076: q = 3'b111;
	13'd1077: q = 3'b111;
	13'd1078: q = 3'b111;
	13'd1079: q = 3'b111;
	13'd1080: q = 3'b111;
	13'd1081: q = 3'b111;
	13'd1082: q = 3'b111;
	13'd1083: q = 3'b111;
	13'd1084: q = 3'b111;
	13'd1085: q = 3'b111;
	13'd1086: q = 3'b000;
	13'd1087: q = 3'b000;
	13'd1088: q = 3'b111;
	13'd1089: q = 3'b111;
	13'd1090: q = 3'b011;
	13'd1091: q = 3'b011;
	13'd1092: q = 3'b011;
	13'd1093: q = 3'b011;
	13'd1094: q = 3'b011;
	13'd1095: q = 3'b011;
	13'd1096: q = 3'b011;
	13'd1097: q = 3'b011;
	13'd1098: q = 3'b011;
	13'd1099: q = 3'b011;
	13'd1100: q = 3'b011;
	13'd1101: q = 3'b011;
	13'd1102: q = 3'b011;
	13'd1103: q = 3'b011;
	13'd1104: q = 3'b011;
	13'd1105: q = 3'b011;
	13'd1106: q = 3'b011;
	13'd1107: q = 3'b011;
	13'd1108: q = 3'b011;
	13'd1109: q = 3'b011;
	13'd1110: q = 3'b011;
	13'd1111: q = 3'b011;
	13'd1112: q = 3'b011;
	13'd1113: q = 3'b011;
	13'd1114: q = 3'b011;
	13'd1115: q = 3'b011;
	13'd1116: q = 3'b011;
	13'd1117: q = 3'b011;
	13'd1118: q = 3'b000;
	13'd1119: q = 3'b000;
	13'd1120: q = 3'b111;
	13'd1121: q = 3'b111;
	13'd1122: q = 3'b011;
	13'd1123: q = 3'b011;
	13'd1124: q = 3'b011;
	13'd1125: q = 3'b011;
	13'd1126: q = 3'b011;
	13'd1127: q = 3'b011;
	13'd1128: q = 3'b011;
	13'd1129: q = 3'b011;
	13'd1130: q = 3'b011;
	13'd1131: q = 3'b011;
	13'd1132: q = 3'b011;
	13'd1133: q = 3'b011;
	13'd1134: q = 3'b011;
	13'd1135: q = 3'b011;
	13'd1136: q = 3'b011;
	13'd1137: q = 3'b011;
	13'd1138: q = 3'b011;
	13'd1139: q = 3'b011;
	13'd1140: q = 3'b011;
	13'd1141: q = 3'b011;
	13'd1142: q = 3'b011;
	13'd1143: q = 3'b011;
	13'd1144: q = 3'b011;
	13'd1145: q = 3'b011;
	13'd1146: q = 3'b011;
	13'd1147: q = 3'b011;
	13'd1148: q = 3'b011;
	13'd1149: q = 3'b011;
	13'd1150: q = 3'b000;
	13'd1151: q = 3'b000;
	13'd1152: q = 3'b111;
	13'd1153: q = 3'b111;
	13'd1154: q = 3'b011;
	13'd1155: q = 3'b011;
	13'd1156: q = 3'b011;
	13'd1157: q = 3'b011;
	13'd1158: q = 3'b011;
	13'd1159: q = 3'b011;
	13'd1160: q = 3'b011;
	13'd1161: q = 3'b011;
	13'd1162: q = 3'b011;
	13'd1163: q = 3'b011;
	13'd1164: q = 3'b011;
	13'd1165: q = 3'b011;
	13'd1166: q = 3'b011;
	13'd1167: q = 3'b011;
	13'd1168: q = 3'b011;
	13'd1169: q = 3'b011;
	13'd1170: q = 3'b011;
	13'd1171: q = 3'b011;
	13'd1172: q = 3'b011;
	13'd1173: q = 3'b011;
	13'd1174: q = 3'b011;
	13'd1175: q = 3'b011;
	13'd1176: q = 3'b011;
	13'd1177: q = 3'b011;
	13'd1178: q = 3'b011;
	13'd1179: q = 3'b011;
	13'd1180: q = 3'b011;
	13'd1181: q = 3'b011;
	13'd1182: q = 3'b000;
	13'd1183: q = 3'b000;
	13'd1184: q = 3'b111;
	13'd1185: q = 3'b111;
	13'd1186: q = 3'b011;
	13'd1187: q = 3'b011;
	13'd1188: q = 3'b011;
	13'd1189: q = 3'b011;
	13'd1190: q = 3'b011;
	13'd1191: q = 3'b011;
	13'd1192: q = 3'b011;
	13'd1193: q = 3'b011;
	13'd1194: q = 3'b011;
	13'd1195: q = 3'b011;
	13'd1196: q = 3'b011;
	13'd1197: q = 3'b011;
	13'd1198: q = 3'b011;
	13'd1199: q = 3'b011;
	13'd1200: q = 3'b011;
	13'd1201: q = 3'b011;
	13'd1202: q = 3'b011;
	13'd1203: q = 3'b011;
	13'd1204: q = 3'b011;
	13'd1205: q = 3'b011;
	13'd1206: q = 3'b011;
	13'd1207: q = 3'b011;
	13'd1208: q = 3'b011;
	13'd1209: q = 3'b011;
	13'd1210: q = 3'b011;
	13'd1211: q = 3'b011;
	13'd1212: q = 3'b011;
	13'd1213: q = 3'b011;
	13'd1214: q = 3'b000;
	13'd1215: q = 3'b000;
	13'd1216: q = 3'b111;
	13'd1217: q = 3'b111;
	13'd1218: q = 3'b011;
	13'd1219: q = 3'b011;
	13'd1220: q = 3'b011;
	13'd1221: q = 3'b011;
	13'd1222: q = 3'b011;
	13'd1223: q = 3'b011;
	13'd1224: q = 3'b011;
	13'd1225: q = 3'b011;
	13'd1226: q = 3'b011;
	13'd1227: q = 3'b011;
	13'd1228: q = 3'b011;
	13'd1229: q = 3'b011;
	13'd1230: q = 3'b011;
	13'd1231: q = 3'b011;
	13'd1232: q = 3'b011;
	13'd1233: q = 3'b011;
	13'd1234: q = 3'b011;
	13'd1235: q = 3'b011;
	13'd1236: q = 3'b011;
	13'd1237: q = 3'b011;
	13'd1238: q = 3'b011;
	13'd1239: q = 3'b011;
	13'd1240: q = 3'b011;
	13'd1241: q = 3'b011;
	13'd1242: q = 3'b011;
	13'd1243: q = 3'b011;
	13'd1244: q = 3'b011;
	13'd1245: q = 3'b011;
	13'd1246: q = 3'b000;
	13'd1247: q = 3'b000;
	13'd1248: q = 3'b111;
	13'd1249: q = 3'b111;
	13'd1250: q = 3'b011;
	13'd1251: q = 3'b011;
	13'd1252: q = 3'b011;
	13'd1253: q = 3'b011;
	13'd1254: q = 3'b011;
	13'd1255: q = 3'b011;
	13'd1256: q = 3'b011;
	13'd1257: q = 3'b011;
	13'd1258: q = 3'b011;
	13'd1259: q = 3'b011;
	13'd1260: q = 3'b011;
	13'd1261: q = 3'b011;
	13'd1262: q = 3'b011;
	13'd1263: q = 3'b011;
	13'd1264: q = 3'b011;
	13'd1265: q = 3'b011;
	13'd1266: q = 3'b011;
	13'd1267: q = 3'b011;
	13'd1268: q = 3'b011;
	13'd1269: q = 3'b011;
	13'd1270: q = 3'b011;
	13'd1271: q = 3'b011;
	13'd1272: q = 3'b011;
	13'd1273: q = 3'b011;
	13'd1274: q = 3'b011;
	13'd1275: q = 3'b011;
	13'd1276: q = 3'b011;
	13'd1277: q = 3'b011;
	13'd1278: q = 3'b000;
	13'd1279: q = 3'b000;
	13'd1280: q = 3'b111;
	13'd1281: q = 3'b111;
	13'd1282: q = 3'b011;
	13'd1283: q = 3'b011;
	13'd1284: q = 3'b011;
	13'd1285: q = 3'b011;
	13'd1286: q = 3'b011;
	13'd1287: q = 3'b011;
	13'd1288: q = 3'b011;
	13'd1289: q = 3'b011;
	13'd1290: q = 3'b011;
	13'd1291: q = 3'b011;
	13'd1292: q = 3'b011;
	13'd1293: q = 3'b011;
	13'd1294: q = 3'b011;
	13'd1295: q = 3'b011;
	13'd1296: q = 3'b011;
	13'd1297: q = 3'b011;
	13'd1298: q = 3'b011;
	13'd1299: q = 3'b011;
	13'd1300: q = 3'b011;
	13'd1301: q = 3'b011;
	13'd1302: q = 3'b011;
	13'd1303: q = 3'b011;
	13'd1304: q = 3'b011;
	13'd1305: q = 3'b011;
	13'd1306: q = 3'b011;
	13'd1307: q = 3'b011;
	13'd1308: q = 3'b011;
	13'd1309: q = 3'b011;
	13'd1310: q = 3'b000;
	13'd1311: q = 3'b000;
	13'd1312: q = 3'b111;
	13'd1313: q = 3'b111;
	13'd1314: q = 3'b011;
	13'd1315: q = 3'b011;
	13'd1316: q = 3'b011;
	13'd1317: q = 3'b011;
	13'd1318: q = 3'b011;
	13'd1319: q = 3'b011;
	13'd1320: q = 3'b011;
	13'd1321: q = 3'b011;
	13'd1322: q = 3'b011;
	13'd1323: q = 3'b011;
	13'd1324: q = 3'b011;
	13'd1325: q = 3'b011;
	13'd1326: q = 3'b011;
	13'd1327: q = 3'b011;
	13'd1328: q = 3'b011;
	13'd1329: q = 3'b011;
	13'd1330: q = 3'b011;
	13'd1331: q = 3'b011;
	13'd1332: q = 3'b011;
	13'd1333: q = 3'b011;
	13'd1334: q = 3'b011;
	13'd1335: q = 3'b011;
	13'd1336: q = 3'b011;
	13'd1337: q = 3'b011;
	13'd1338: q = 3'b011;
	13'd1339: q = 3'b011;
	13'd1340: q = 3'b011;
	13'd1341: q = 3'b011;
	13'd1342: q = 3'b000;
	13'd1343: q = 3'b000;
	13'd1344: q = 3'b111;
	13'd1345: q = 3'b111;
	13'd1346: q = 3'b011;
	13'd1347: q = 3'b011;
	13'd1348: q = 3'b011;
	13'd1349: q = 3'b011;
	13'd1350: q = 3'b011;
	13'd1351: q = 3'b011;
	13'd1352: q = 3'b011;
	13'd1353: q = 3'b011;
	13'd1354: q = 3'b011;
	13'd1355: q = 3'b011;
	13'd1356: q = 3'b011;
	13'd1357: q = 3'b011;
	13'd1358: q = 3'b011;
	13'd1359: q = 3'b011;
	13'd1360: q = 3'b011;
	13'd1361: q = 3'b011;
	13'd1362: q = 3'b011;
	13'd1363: q = 3'b011;
	13'd1364: q = 3'b011;
	13'd1365: q = 3'b011;
	13'd1366: q = 3'b011;
	13'd1367: q = 3'b011;
	13'd1368: q = 3'b011;
	13'd1369: q = 3'b011;
	13'd1370: q = 3'b011;
	13'd1371: q = 3'b011;
	13'd1372: q = 3'b011;
	13'd1373: q = 3'b011;
	13'd1374: q = 3'b000;
	13'd1375: q = 3'b000;
	13'd1376: q = 3'b111;
	13'd1377: q = 3'b111;
	13'd1378: q = 3'b011;
	13'd1379: q = 3'b011;
	13'd1380: q = 3'b011;
	13'd1381: q = 3'b011;
	13'd1382: q = 3'b011;
	13'd1383: q = 3'b011;
	13'd1384: q = 3'b011;
	13'd1385: q = 3'b011;
	13'd1386: q = 3'b011;
	13'd1387: q = 3'b011;
	13'd1388: q = 3'b011;
	13'd1389: q = 3'b011;
	13'd1390: q = 3'b011;
	13'd1391: q = 3'b011;
	13'd1392: q = 3'b011;
	13'd1393: q = 3'b011;
	13'd1394: q = 3'b011;
	13'd1395: q = 3'b011;
	13'd1396: q = 3'b011;
	13'd1397: q = 3'b011;
	13'd1398: q = 3'b011;
	13'd1399: q = 3'b011;
	13'd1400: q = 3'b011;
	13'd1401: q = 3'b011;
	13'd1402: q = 3'b011;
	13'd1403: q = 3'b011;
	13'd1404: q = 3'b011;
	13'd1405: q = 3'b011;
	13'd1406: q = 3'b000;
	13'd1407: q = 3'b000;
	13'd1408: q = 3'b111;
	13'd1409: q = 3'b111;
	13'd1410: q = 3'b011;
	13'd1411: q = 3'b011;
	13'd1412: q = 3'b011;
	13'd1413: q = 3'b011;
	13'd1414: q = 3'b011;
	13'd1415: q = 3'b011;
	13'd1416: q = 3'b011;
	13'd1417: q = 3'b011;
	13'd1418: q = 3'b011;
	13'd1419: q = 3'b011;
	13'd1420: q = 3'b011;
	13'd1421: q = 3'b011;
	13'd1422: q = 3'b011;
	13'd1423: q = 3'b011;
	13'd1424: q = 3'b011;
	13'd1425: q = 3'b011;
	13'd1426: q = 3'b011;
	13'd1427: q = 3'b011;
	13'd1428: q = 3'b011;
	13'd1429: q = 3'b011;
	13'd1430: q = 3'b011;
	13'd1431: q = 3'b011;
	13'd1432: q = 3'b011;
	13'd1433: q = 3'b011;
	13'd1434: q = 3'b011;
	13'd1435: q = 3'b011;
	13'd1436: q = 3'b011;
	13'd1437: q = 3'b011;
	13'd1438: q = 3'b000;
	13'd1439: q = 3'b000;
	13'd1440: q = 3'b111;
	13'd1441: q = 3'b111;
	13'd1442: q = 3'b011;
	13'd1443: q = 3'b011;
	13'd1444: q = 3'b011;
	13'd1445: q = 3'b011;
	13'd1446: q = 3'b011;
	13'd1447: q = 3'b011;
	13'd1448: q = 3'b011;
	13'd1449: q = 3'b011;
	13'd1450: q = 3'b011;
	13'd1451: q = 3'b011;
	13'd1452: q = 3'b011;
	13'd1453: q = 3'b011;
	13'd1454: q = 3'b011;
	13'd1455: q = 3'b011;
	13'd1456: q = 3'b011;
	13'd1457: q = 3'b011;
	13'd1458: q = 3'b011;
	13'd1459: q = 3'b011;
	13'd1460: q = 3'b011;
	13'd1461: q = 3'b011;
	13'd1462: q = 3'b011;
	13'd1463: q = 3'b011;
	13'd1464: q = 3'b011;
	13'd1465: q = 3'b011;
	13'd1466: q = 3'b011;
	13'd1467: q = 3'b011;
	13'd1468: q = 3'b011;
	13'd1469: q = 3'b011;
	13'd1470: q = 3'b000;
	13'd1471: q = 3'b000;
	13'd1472: q = 3'b111;
	13'd1473: q = 3'b111;
	13'd1474: q = 3'b011;
	13'd1475: q = 3'b011;
	13'd1476: q = 3'b011;
	13'd1477: q = 3'b011;
	13'd1478: q = 3'b011;
	13'd1479: q = 3'b011;
	13'd1480: q = 3'b011;
	13'd1481: q = 3'b011;
	13'd1482: q = 3'b011;
	13'd1483: q = 3'b011;
	13'd1484: q = 3'b011;
	13'd1485: q = 3'b011;
	13'd1486: q = 3'b011;
	13'd1487: q = 3'b011;
	13'd1488: q = 3'b011;
	13'd1489: q = 3'b011;
	13'd1490: q = 3'b011;
	13'd1491: q = 3'b011;
	13'd1492: q = 3'b011;
	13'd1493: q = 3'b011;
	13'd1494: q = 3'b011;
	13'd1495: q = 3'b011;
	13'd1496: q = 3'b011;
	13'd1497: q = 3'b011;
	13'd1498: q = 3'b011;
	13'd1499: q = 3'b011;
	13'd1500: q = 3'b011;
	13'd1501: q = 3'b011;
	13'd1502: q = 3'b000;
	13'd1503: q = 3'b000;
	13'd1504: q = 3'b111;
	13'd1505: q = 3'b111;
	13'd1506: q = 3'b011;
	13'd1507: q = 3'b011;
	13'd1508: q = 3'b011;
	13'd1509: q = 3'b011;
	13'd1510: q = 3'b011;
	13'd1511: q = 3'b011;
	13'd1512: q = 3'b011;
	13'd1513: q = 3'b011;
	13'd1514: q = 3'b011;
	13'd1515: q = 3'b011;
	13'd1516: q = 3'b011;
	13'd1517: q = 3'b011;
	13'd1518: q = 3'b011;
	13'd1519: q = 3'b011;
	13'd1520: q = 3'b011;
	13'd1521: q = 3'b011;
	13'd1522: q = 3'b011;
	13'd1523: q = 3'b011;
	13'd1524: q = 3'b011;
	13'd1525: q = 3'b011;
	13'd1526: q = 3'b011;
	13'd1527: q = 3'b011;
	13'd1528: q = 3'b011;
	13'd1529: q = 3'b011;
	13'd1530: q = 3'b011;
	13'd1531: q = 3'b011;
	13'd1532: q = 3'b011;
	13'd1533: q = 3'b011;
	13'd1534: q = 3'b000;
	13'd1535: q = 3'b000;
	13'd1536: q = 3'b111;
	13'd1537: q = 3'b111;
	13'd1538: q = 3'b011;
	13'd1539: q = 3'b011;
	13'd1540: q = 3'b011;
	13'd1541: q = 3'b011;
	13'd1542: q = 3'b011;
	13'd1543: q = 3'b011;
	13'd1544: q = 3'b011;
	13'd1545: q = 3'b011;
	13'd1546: q = 3'b011;
	13'd1547: q = 3'b011;
	13'd1548: q = 3'b011;
	13'd1549: q = 3'b011;
	13'd1550: q = 3'b011;
	13'd1551: q = 3'b011;
	13'd1552: q = 3'b011;
	13'd1553: q = 3'b011;
	13'd1554: q = 3'b011;
	13'd1555: q = 3'b011;
	13'd1556: q = 3'b011;
	13'd1557: q = 3'b011;
	13'd1558: q = 3'b011;
	13'd1559: q = 3'b011;
	13'd1560: q = 3'b011;
	13'd1561: q = 3'b011;
	13'd1562: q = 3'b011;
	13'd1563: q = 3'b011;
	13'd1564: q = 3'b011;
	13'd1565: q = 3'b011;
	13'd1566: q = 3'b000;
	13'd1567: q = 3'b000;
	13'd1568: q = 3'b111;
	13'd1569: q = 3'b111;
	13'd1570: q = 3'b011;
	13'd1571: q = 3'b011;
	13'd1572: q = 3'b011;
	13'd1573: q = 3'b011;
	13'd1574: q = 3'b011;
	13'd1575: q = 3'b011;
	13'd1576: q = 3'b011;
	13'd1577: q = 3'b011;
	13'd1578: q = 3'b011;
	13'd1579: q = 3'b011;
	13'd1580: q = 3'b011;
	13'd1581: q = 3'b011;
	13'd1582: q = 3'b011;
	13'd1583: q = 3'b011;
	13'd1584: q = 3'b011;
	13'd1585: q = 3'b011;
	13'd1586: q = 3'b011;
	13'd1587: q = 3'b011;
	13'd1588: q = 3'b011;
	13'd1589: q = 3'b011;
	13'd1590: q = 3'b011;
	13'd1591: q = 3'b011;
	13'd1592: q = 3'b011;
	13'd1593: q = 3'b011;
	13'd1594: q = 3'b011;
	13'd1595: q = 3'b011;
	13'd1596: q = 3'b011;
	13'd1597: q = 3'b011;
	13'd1598: q = 3'b000;
	13'd1599: q = 3'b000;
	13'd1600: q = 3'b111;
	13'd1601: q = 3'b111;
	13'd1602: q = 3'b011;
	13'd1603: q = 3'b011;
	13'd1604: q = 3'b011;
	13'd1605: q = 3'b011;
	13'd1606: q = 3'b011;
	13'd1607: q = 3'b011;
	13'd1608: q = 3'b011;
	13'd1609: q = 3'b011;
	13'd1610: q = 3'b011;
	13'd1611: q = 3'b011;
	13'd1612: q = 3'b011;
	13'd1613: q = 3'b011;
	13'd1614: q = 3'b011;
	13'd1615: q = 3'b011;
	13'd1616: q = 3'b011;
	13'd1617: q = 3'b011;
	13'd1618: q = 3'b011;
	13'd1619: q = 3'b011;
	13'd1620: q = 3'b011;
	13'd1621: q = 3'b011;
	13'd1622: q = 3'b011;
	13'd1623: q = 3'b011;
	13'd1624: q = 3'b011;
	13'd1625: q = 3'b011;
	13'd1626: q = 3'b011;
	13'd1627: q = 3'b011;
	13'd1628: q = 3'b011;
	13'd1629: q = 3'b011;
	13'd1630: q = 3'b000;
	13'd1631: q = 3'b000;
	13'd1632: q = 3'b111;
	13'd1633: q = 3'b111;
	13'd1634: q = 3'b011;
	13'd1635: q = 3'b011;
	13'd1636: q = 3'b011;
	13'd1637: q = 3'b011;
	13'd1638: q = 3'b011;
	13'd1639: q = 3'b011;
	13'd1640: q = 3'b011;
	13'd1641: q = 3'b011;
	13'd1642: q = 3'b011;
	13'd1643: q = 3'b011;
	13'd1644: q = 3'b011;
	13'd1645: q = 3'b011;
	13'd1646: q = 3'b011;
	13'd1647: q = 3'b011;
	13'd1648: q = 3'b011;
	13'd1649: q = 3'b011;
	13'd1650: q = 3'b011;
	13'd1651: q = 3'b011;
	13'd1652: q = 3'b011;
	13'd1653: q = 3'b011;
	13'd1654: q = 3'b011;
	13'd1655: q = 3'b011;
	13'd1656: q = 3'b011;
	13'd1657: q = 3'b011;
	13'd1658: q = 3'b011;
	13'd1659: q = 3'b011;
	13'd1660: q = 3'b011;
	13'd1661: q = 3'b011;
	13'd1662: q = 3'b000;
	13'd1663: q = 3'b000;
	13'd1664: q = 3'b111;
	13'd1665: q = 3'b111;
	13'd1666: q = 3'b011;
	13'd1667: q = 3'b011;
	13'd1668: q = 3'b011;
	13'd1669: q = 3'b011;
	13'd1670: q = 3'b011;
	13'd1671: q = 3'b011;
	13'd1672: q = 3'b011;
	13'd1673: q = 3'b011;
	13'd1674: q = 3'b011;
	13'd1675: q = 3'b011;
	13'd1676: q = 3'b011;
	13'd1677: q = 3'b011;
	13'd1678: q = 3'b011;
	13'd1679: q = 3'b011;
	13'd1680: q = 3'b011;
	13'd1681: q = 3'b011;
	13'd1682: q = 3'b011;
	13'd1683: q = 3'b011;
	13'd1684: q = 3'b011;
	13'd1685: q = 3'b011;
	13'd1686: q = 3'b011;
	13'd1687: q = 3'b011;
	13'd1688: q = 3'b011;
	13'd1689: q = 3'b011;
	13'd1690: q = 3'b011;
	13'd1691: q = 3'b011;
	13'd1692: q = 3'b011;
	13'd1693: q = 3'b011;
	13'd1694: q = 3'b000;
	13'd1695: q = 3'b000;
	13'd1696: q = 3'b111;
	13'd1697: q = 3'b111;
	13'd1698: q = 3'b011;
	13'd1699: q = 3'b011;
	13'd1700: q = 3'b011;
	13'd1701: q = 3'b011;
	13'd1702: q = 3'b011;
	13'd1703: q = 3'b011;
	13'd1704: q = 3'b011;
	13'd1705: q = 3'b011;
	13'd1706: q = 3'b011;
	13'd1707: q = 3'b011;
	13'd1708: q = 3'b011;
	13'd1709: q = 3'b011;
	13'd1710: q = 3'b011;
	13'd1711: q = 3'b011;
	13'd1712: q = 3'b011;
	13'd1713: q = 3'b011;
	13'd1714: q = 3'b011;
	13'd1715: q = 3'b011;
	13'd1716: q = 3'b011;
	13'd1717: q = 3'b011;
	13'd1718: q = 3'b011;
	13'd1719: q = 3'b011;
	13'd1720: q = 3'b011;
	13'd1721: q = 3'b011;
	13'd1722: q = 3'b011;
	13'd1723: q = 3'b011;
	13'd1724: q = 3'b011;
	13'd1725: q = 3'b011;
	13'd1726: q = 3'b000;
	13'd1727: q = 3'b000;
	13'd1728: q = 3'b111;
	13'd1729: q = 3'b111;
	13'd1730: q = 3'b011;
	13'd1731: q = 3'b011;
	13'd1732: q = 3'b011;
	13'd1733: q = 3'b011;
	13'd1734: q = 3'b011;
	13'd1735: q = 3'b011;
	13'd1736: q = 3'b011;
	13'd1737: q = 3'b011;
	13'd1738: q = 3'b011;
	13'd1739: q = 3'b011;
	13'd1740: q = 3'b011;
	13'd1741: q = 3'b011;
	13'd1742: q = 3'b011;
	13'd1743: q = 3'b011;
	13'd1744: q = 3'b011;
	13'd1745: q = 3'b011;
	13'd1746: q = 3'b011;
	13'd1747: q = 3'b011;
	13'd1748: q = 3'b011;
	13'd1749: q = 3'b011;
	13'd1750: q = 3'b011;
	13'd1751: q = 3'b011;
	13'd1752: q = 3'b011;
	13'd1753: q = 3'b011;
	13'd1754: q = 3'b011;
	13'd1755: q = 3'b011;
	13'd1756: q = 3'b011;
	13'd1757: q = 3'b011;
	13'd1758: q = 3'b000;
	13'd1759: q = 3'b000;
	13'd1760: q = 3'b111;
	13'd1761: q = 3'b111;
	13'd1762: q = 3'b011;
	13'd1763: q = 3'b011;
	13'd1764: q = 3'b011;
	13'd1765: q = 3'b011;
	13'd1766: q = 3'b011;
	13'd1767: q = 3'b011;
	13'd1768: q = 3'b011;
	13'd1769: q = 3'b011;
	13'd1770: q = 3'b011;
	13'd1771: q = 3'b011;
	13'd1772: q = 3'b011;
	13'd1773: q = 3'b011;
	13'd1774: q = 3'b011;
	13'd1775: q = 3'b011;
	13'd1776: q = 3'b011;
	13'd1777: q = 3'b011;
	13'd1778: q = 3'b011;
	13'd1779: q = 3'b011;
	13'd1780: q = 3'b011;
	13'd1781: q = 3'b011;
	13'd1782: q = 3'b011;
	13'd1783: q = 3'b011;
	13'd1784: q = 3'b011;
	13'd1785: q = 3'b011;
	13'd1786: q = 3'b011;
	13'd1787: q = 3'b011;
	13'd1788: q = 3'b011;
	13'd1789: q = 3'b011;
	13'd1790: q = 3'b000;
	13'd1791: q = 3'b000;
	13'd1792: q = 3'b111;
	13'd1793: q = 3'b111;
	13'd1794: q = 3'b011;
	13'd1795: q = 3'b011;
	13'd1796: q = 3'b011;
	13'd1797: q = 3'b011;
	13'd1798: q = 3'b011;
	13'd1799: q = 3'b011;
	13'd1800: q = 3'b011;
	13'd1801: q = 3'b011;
	13'd1802: q = 3'b011;
	13'd1803: q = 3'b011;
	13'd1804: q = 3'b011;
	13'd1805: q = 3'b011;
	13'd1806: q = 3'b011;
	13'd1807: q = 3'b011;
	13'd1808: q = 3'b011;
	13'd1809: q = 3'b011;
	13'd1810: q = 3'b011;
	13'd1811: q = 3'b011;
	13'd1812: q = 3'b011;
	13'd1813: q = 3'b011;
	13'd1814: q = 3'b011;
	13'd1815: q = 3'b011;
	13'd1816: q = 3'b011;
	13'd1817: q = 3'b011;
	13'd1818: q = 3'b011;
	13'd1819: q = 3'b011;
	13'd1820: q = 3'b011;
	13'd1821: q = 3'b011;
	13'd1822: q = 3'b000;
	13'd1823: q = 3'b000;
	13'd1824: q = 3'b111;
	13'd1825: q = 3'b111;
	13'd1826: q = 3'b011;
	13'd1827: q = 3'b011;
	13'd1828: q = 3'b011;
	13'd1829: q = 3'b011;
	13'd1830: q = 3'b011;
	13'd1831: q = 3'b011;
	13'd1832: q = 3'b011;
	13'd1833: q = 3'b011;
	13'd1834: q = 3'b011;
	13'd1835: q = 3'b011;
	13'd1836: q = 3'b011;
	13'd1837: q = 3'b011;
	13'd1838: q = 3'b011;
	13'd1839: q = 3'b011;
	13'd1840: q = 3'b011;
	13'd1841: q = 3'b011;
	13'd1842: q = 3'b011;
	13'd1843: q = 3'b011;
	13'd1844: q = 3'b011;
	13'd1845: q = 3'b011;
	13'd1846: q = 3'b011;
	13'd1847: q = 3'b011;
	13'd1848: q = 3'b011;
	13'd1849: q = 3'b011;
	13'd1850: q = 3'b011;
	13'd1851: q = 3'b011;
	13'd1852: q = 3'b011;
	13'd1853: q = 3'b011;
	13'd1854: q = 3'b000;
	13'd1855: q = 3'b000;
	13'd1856: q = 3'b111;
	13'd1857: q = 3'b111;
	13'd1858: q = 3'b011;
	13'd1859: q = 3'b011;
	13'd1860: q = 3'b011;
	13'd1861: q = 3'b011;
	13'd1862: q = 3'b011;
	13'd1863: q = 3'b011;
	13'd1864: q = 3'b011;
	13'd1865: q = 3'b011;
	13'd1866: q = 3'b011;
	13'd1867: q = 3'b011;
	13'd1868: q = 3'b011;
	13'd1869: q = 3'b011;
	13'd1870: q = 3'b011;
	13'd1871: q = 3'b011;
	13'd1872: q = 3'b011;
	13'd1873: q = 3'b011;
	13'd1874: q = 3'b011;
	13'd1875: q = 3'b011;
	13'd1876: q = 3'b011;
	13'd1877: q = 3'b011;
	13'd1878: q = 3'b011;
	13'd1879: q = 3'b011;
	13'd1880: q = 3'b011;
	13'd1881: q = 3'b011;
	13'd1882: q = 3'b011;
	13'd1883: q = 3'b011;
	13'd1884: q = 3'b011;
	13'd1885: q = 3'b011;
	13'd1886: q = 3'b000;
	13'd1887: q = 3'b000;
	13'd1888: q = 3'b111;
	13'd1889: q = 3'b111;
	13'd1890: q = 3'b011;
	13'd1891: q = 3'b011;
	13'd1892: q = 3'b011;
	13'd1893: q = 3'b011;
	13'd1894: q = 3'b011;
	13'd1895: q = 3'b011;
	13'd1896: q = 3'b011;
	13'd1897: q = 3'b011;
	13'd1898: q = 3'b011;
	13'd1899: q = 3'b011;
	13'd1900: q = 3'b011;
	13'd1901: q = 3'b011;
	13'd1902: q = 3'b011;
	13'd1903: q = 3'b011;
	13'd1904: q = 3'b011;
	13'd1905: q = 3'b011;
	13'd1906: q = 3'b011;
	13'd1907: q = 3'b011;
	13'd1908: q = 3'b011;
	13'd1909: q = 3'b011;
	13'd1910: q = 3'b011;
	13'd1911: q = 3'b011;
	13'd1912: q = 3'b011;
	13'd1913: q = 3'b011;
	13'd1914: q = 3'b011;
	13'd1915: q = 3'b011;
	13'd1916: q = 3'b011;
	13'd1917: q = 3'b011;
	13'd1918: q = 3'b000;
	13'd1919: q = 3'b000;
	13'd1920: q = 3'b111;
	13'd1921: q = 3'b111;
	13'd1922: q = 3'b011;
	13'd1923: q = 3'b011;
	13'd1924: q = 3'b011;
	13'd1925: q = 3'b011;
	13'd1926: q = 3'b011;
	13'd1927: q = 3'b011;
	13'd1928: q = 3'b011;
	13'd1929: q = 3'b011;
	13'd1930: q = 3'b011;
	13'd1931: q = 3'b011;
	13'd1932: q = 3'b011;
	13'd1933: q = 3'b011;
	13'd1934: q = 3'b011;
	13'd1935: q = 3'b011;
	13'd1936: q = 3'b011;
	13'd1937: q = 3'b011;
	13'd1938: q = 3'b011;
	13'd1939: q = 3'b011;
	13'd1940: q = 3'b011;
	13'd1941: q = 3'b011;
	13'd1942: q = 3'b011;
	13'd1943: q = 3'b011;
	13'd1944: q = 3'b011;
	13'd1945: q = 3'b011;
	13'd1946: q = 3'b011;
	13'd1947: q = 3'b011;
	13'd1948: q = 3'b011;
	13'd1949: q = 3'b011;
	13'd1950: q = 3'b000;
	13'd1951: q = 3'b000;
	13'd1952: q = 3'b111;
	13'd1953: q = 3'b111;
	13'd1954: q = 3'b011;
	13'd1955: q = 3'b011;
	13'd1956: q = 3'b011;
	13'd1957: q = 3'b011;
	13'd1958: q = 3'b011;
	13'd1959: q = 3'b011;
	13'd1960: q = 3'b011;
	13'd1961: q = 3'b011;
	13'd1962: q = 3'b011;
	13'd1963: q = 3'b011;
	13'd1964: q = 3'b011;
	13'd1965: q = 3'b011;
	13'd1966: q = 3'b011;
	13'd1967: q = 3'b011;
	13'd1968: q = 3'b011;
	13'd1969: q = 3'b011;
	13'd1970: q = 3'b011;
	13'd1971: q = 3'b011;
	13'd1972: q = 3'b011;
	13'd1973: q = 3'b011;
	13'd1974: q = 3'b011;
	13'd1975: q = 3'b011;
	13'd1976: q = 3'b011;
	13'd1977: q = 3'b011;
	13'd1978: q = 3'b011;
	13'd1979: q = 3'b011;
	13'd1980: q = 3'b011;
	13'd1981: q = 3'b011;
	13'd1982: q = 3'b000;
	13'd1983: q = 3'b000;
	13'd1984: q = 3'b000;
	13'd1985: q = 3'b000;
	13'd1986: q = 3'b000;
	13'd1987: q = 3'b000;
	13'd1988: q = 3'b000;
	13'd1989: q = 3'b000;
	13'd1990: q = 3'b000;
	13'd1991: q = 3'b000;
	13'd1992: q = 3'b000;
	13'd1993: q = 3'b000;
	13'd1994: q = 3'b000;
	13'd1995: q = 3'b000;
	13'd1996: q = 3'b000;
	13'd1997: q = 3'b000;
	13'd1998: q = 3'b000;
	13'd1999: q = 3'b000;
	13'd2000: q = 3'b000;
	13'd2001: q = 3'b000;
	13'd2002: q = 3'b000;
	13'd2003: q = 3'b000;
	13'd2004: q = 3'b000;
	13'd2005: q = 3'b000;
	13'd2006: q = 3'b000;
	13'd2007: q = 3'b000;
	13'd2008: q = 3'b000;
	13'd2009: q = 3'b000;
	13'd2010: q = 3'b000;
	13'd2011: q = 3'b000;
	13'd2012: q = 3'b000;
	13'd2013: q = 3'b000;
	13'd2014: q = 3'b000;
	13'd2015: q = 3'b000;
	13'd2016: q = 3'b000;
	13'd2017: q = 3'b000;
	13'd2018: q = 3'b000;
	13'd2019: q = 3'b000;
	13'd2020: q = 3'b000;
	13'd2021: q = 3'b000;
	13'd2022: q = 3'b000;
	13'd2023: q = 3'b000;
	13'd2024: q = 3'b000;
	13'd2025: q = 3'b000;
	13'd2026: q = 3'b000;
	13'd2027: q = 3'b000;
	13'd2028: q = 3'b000;
	13'd2029: q = 3'b000;
	13'd2030: q = 3'b000;
	13'd2031: q = 3'b000;
	13'd2032: q = 3'b000;
	13'd2033: q = 3'b000;
	13'd2034: q = 3'b000;
	13'd2035: q = 3'b000;
	13'd2036: q = 3'b000;
	13'd2037: q = 3'b000;
	13'd2038: q = 3'b000;
	13'd2039: q = 3'b000;
	13'd2040: q = 3'b000;
	13'd2041: q = 3'b000;
	13'd2042: q = 3'b000;
	13'd2043: q = 3'b000;
	13'd2044: q = 3'b000;
	13'd2045: q = 3'b000;
	13'd2046: q = 3'b000;
	13'd2047: q = 3'b000;
	13'd2048: q = 3'b000;
	13'd2049: q = 3'b000;
	13'd2050: q = 3'b000;
	13'd2051: q = 3'b000;
	13'd2052: q = 3'b000;
	13'd2053: q = 3'b000;
	13'd2054: q = 3'b000;
	13'd2055: q = 3'b000;
	13'd2056: q = 3'b000;
	13'd2057: q = 3'b000;
	13'd2058: q = 3'b000;
	13'd2059: q = 3'b000;
	13'd2060: q = 3'b000;
	13'd2061: q = 3'b000;
	13'd2062: q = 3'b000;
	13'd2063: q = 3'b000;
	13'd2064: q = 3'b000;
	13'd2065: q = 3'b000;
	13'd2066: q = 3'b000;
	13'd2067: q = 3'b000;
	13'd2068: q = 3'b000;
	13'd2069: q = 3'b000;
	13'd2070: q = 3'b000;
	13'd2071: q = 3'b000;
	13'd2072: q = 3'b000;
	13'd2073: q = 3'b000;
	13'd2074: q = 3'b000;
	13'd2075: q = 3'b000;
	13'd2076: q = 3'b000;
	13'd2077: q = 3'b000;
	13'd2078: q = 3'b000;
	13'd2079: q = 3'b000;
	13'd2080: q = 3'b000;
	13'd2081: q = 3'b000;
	13'd2082: q = 3'b000;
	13'd2083: q = 3'b000;
	13'd2084: q = 3'b000;
	13'd2085: q = 3'b000;
	13'd2086: q = 3'b000;
	13'd2087: q = 3'b000;
	13'd2088: q = 3'b000;
	13'd2089: q = 3'b000;
	13'd2090: q = 3'b000;
	13'd2091: q = 3'b000;
	13'd2092: q = 3'b000;
	13'd2093: q = 3'b000;
	13'd2094: q = 3'b000;
	13'd2095: q = 3'b000;
	13'd2096: q = 3'b000;
	13'd2097: q = 3'b000;
	13'd2098: q = 3'b000;
	13'd2099: q = 3'b000;
	13'd2100: q = 3'b000;
	13'd2101: q = 3'b000;
	13'd2102: q = 3'b000;
	13'd2103: q = 3'b000;
	13'd2104: q = 3'b000;
	13'd2105: q = 3'b000;
	13'd2106: q = 3'b000;
	13'd2107: q = 3'b000;
	13'd2108: q = 3'b000;
	13'd2109: q = 3'b000;
	13'd2110: q = 3'b000;
	13'd2111: q = 3'b000;
	13'd2112: q = 3'b000;
	13'd2113: q = 3'b000;
	13'd2114: q = 3'b111;
	13'd2115: q = 3'b111;
	13'd2116: q = 3'b111;
	13'd2117: q = 3'b111;
	13'd2118: q = 3'b111;
	13'd2119: q = 3'b111;
	13'd2120: q = 3'b111;
	13'd2121: q = 3'b111;
	13'd2122: q = 3'b111;
	13'd2123: q = 3'b111;
	13'd2124: q = 3'b111;
	13'd2125: q = 3'b111;
	13'd2126: q = 3'b111;
	13'd2127: q = 3'b111;
	13'd2128: q = 3'b111;
	13'd2129: q = 3'b111;
	13'd2130: q = 3'b111;
	13'd2131: q = 3'b111;
	13'd2132: q = 3'b111;
	13'd2133: q = 3'b111;
	13'd2134: q = 3'b111;
	13'd2135: q = 3'b111;
	13'd2136: q = 3'b111;
	13'd2137: q = 3'b111;
	13'd2138: q = 3'b111;
	13'd2139: q = 3'b111;
	13'd2140: q = 3'b111;
	13'd2141: q = 3'b111;
	13'd2142: q = 3'b000;
	13'd2143: q = 3'b000;
	13'd2144: q = 3'b000;
	13'd2145: q = 3'b000;
	13'd2146: q = 3'b111;
	13'd2147: q = 3'b111;
	13'd2148: q = 3'b111;
	13'd2149: q = 3'b111;
	13'd2150: q = 3'b111;
	13'd2151: q = 3'b111;
	13'd2152: q = 3'b111;
	13'd2153: q = 3'b111;
	13'd2154: q = 3'b111;
	13'd2155: q = 3'b111;
	13'd2156: q = 3'b111;
	13'd2157: q = 3'b111;
	13'd2158: q = 3'b111;
	13'd2159: q = 3'b111;
	13'd2160: q = 3'b111;
	13'd2161: q = 3'b111;
	13'd2162: q = 3'b111;
	13'd2163: q = 3'b111;
	13'd2164: q = 3'b111;
	13'd2165: q = 3'b111;
	13'd2166: q = 3'b111;
	13'd2167: q = 3'b111;
	13'd2168: q = 3'b111;
	13'd2169: q = 3'b111;
	13'd2170: q = 3'b111;
	13'd2171: q = 3'b111;
	13'd2172: q = 3'b111;
	13'd2173: q = 3'b111;
	13'd2174: q = 3'b000;
	13'd2175: q = 3'b000;
	13'd2176: q = 3'b111;
	13'd2177: q = 3'b111;
	13'd2178: q = 3'b011;
	13'd2179: q = 3'b011;
	13'd2180: q = 3'b011;
	13'd2181: q = 3'b011;
	13'd2182: q = 3'b011;
	13'd2183: q = 3'b011;
	13'd2184: q = 3'b011;
	13'd2185: q = 3'b011;
	13'd2186: q = 3'b011;
	13'd2187: q = 3'b011;
	13'd2188: q = 3'b011;
	13'd2189: q = 3'b011;
	13'd2190: q = 3'b011;
	13'd2191: q = 3'b011;
	13'd2192: q = 3'b011;
	13'd2193: q = 3'b011;
	13'd2194: q = 3'b011;
	13'd2195: q = 3'b011;
	13'd2196: q = 3'b011;
	13'd2197: q = 3'b011;
	13'd2198: q = 3'b011;
	13'd2199: q = 3'b011;
	13'd2200: q = 3'b011;
	13'd2201: q = 3'b011;
	13'd2202: q = 3'b011;
	13'd2203: q = 3'b011;
	13'd2204: q = 3'b011;
	13'd2205: q = 3'b011;
	13'd2206: q = 3'b000;
	13'd2207: q = 3'b000;
	13'd2208: q = 3'b111;
	13'd2209: q = 3'b111;
	13'd2210: q = 3'b011;
	13'd2211: q = 3'b011;
	13'd2212: q = 3'b011;
	13'd2213: q = 3'b011;
	13'd2214: q = 3'b011;
	13'd2215: q = 3'b011;
	13'd2216: q = 3'b011;
	13'd2217: q = 3'b011;
	13'd2218: q = 3'b011;
	13'd2219: q = 3'b011;
	13'd2220: q = 3'b011;
	13'd2221: q = 3'b011;
	13'd2222: q = 3'b011;
	13'd2223: q = 3'b011;
	13'd2224: q = 3'b011;
	13'd2225: q = 3'b011;
	13'd2226: q = 3'b011;
	13'd2227: q = 3'b011;
	13'd2228: q = 3'b011;
	13'd2229: q = 3'b011;
	13'd2230: q = 3'b011;
	13'd2231: q = 3'b011;
	13'd2232: q = 3'b011;
	13'd2233: q = 3'b011;
	13'd2234: q = 3'b011;
	13'd2235: q = 3'b011;
	13'd2236: q = 3'b011;
	13'd2237: q = 3'b011;
	13'd2238: q = 3'b000;
	13'd2239: q = 3'b000;
	13'd2240: q = 3'b111;
	13'd2241: q = 3'b111;
	13'd2242: q = 3'b011;
	13'd2243: q = 3'b011;
	13'd2244: q = 3'b011;
	13'd2245: q = 3'b011;
	13'd2246: q = 3'b011;
	13'd2247: q = 3'b011;
	13'd2248: q = 3'b011;
	13'd2249: q = 3'b011;
	13'd2250: q = 3'b011;
	13'd2251: q = 3'b011;
	13'd2252: q = 3'b011;
	13'd2253: q = 3'b011;
	13'd2254: q = 3'b011;
	13'd2255: q = 3'b011;
	13'd2256: q = 3'b011;
	13'd2257: q = 3'b011;
	13'd2258: q = 3'b011;
	13'd2259: q = 3'b011;
	13'd2260: q = 3'b011;
	13'd2261: q = 3'b011;
	13'd2262: q = 3'b011;
	13'd2263: q = 3'b011;
	13'd2264: q = 3'b011;
	13'd2265: q = 3'b011;
	13'd2266: q = 3'b011;
	13'd2267: q = 3'b011;
	13'd2268: q = 3'b011;
	13'd2269: q = 3'b011;
	13'd2270: q = 3'b000;
	13'd2271: q = 3'b000;
	13'd2272: q = 3'b111;
	13'd2273: q = 3'b111;
	13'd2274: q = 3'b011;
	13'd2275: q = 3'b011;
	13'd2276: q = 3'b011;
	13'd2277: q = 3'b011;
	13'd2278: q = 3'b011;
	13'd2279: q = 3'b011;
	13'd2280: q = 3'b011;
	13'd2281: q = 3'b011;
	13'd2282: q = 3'b011;
	13'd2283: q = 3'b011;
	13'd2284: q = 3'b011;
	13'd2285: q = 3'b011;
	13'd2286: q = 3'b011;
	13'd2287: q = 3'b011;
	13'd2288: q = 3'b011;
	13'd2289: q = 3'b011;
	13'd2290: q = 3'b011;
	13'd2291: q = 3'b011;
	13'd2292: q = 3'b011;
	13'd2293: q = 3'b011;
	13'd2294: q = 3'b011;
	13'd2295: q = 3'b011;
	13'd2296: q = 3'b011;
	13'd2297: q = 3'b011;
	13'd2298: q = 3'b011;
	13'd2299: q = 3'b011;
	13'd2300: q = 3'b011;
	13'd2301: q = 3'b011;
	13'd2302: q = 3'b000;
	13'd2303: q = 3'b000;
	13'd2304: q = 3'b111;
	13'd2305: q = 3'b111;
	13'd2306: q = 3'b011;
	13'd2307: q = 3'b011;
	13'd2308: q = 3'b011;
	13'd2309: q = 3'b011;
	13'd2310: q = 3'b011;
	13'd2311: q = 3'b011;
	13'd2312: q = 3'b011;
	13'd2313: q = 3'b011;
	13'd2314: q = 3'b011;
	13'd2315: q = 3'b011;
	13'd2316: q = 3'b011;
	13'd2317: q = 3'b011;
	13'd2318: q = 3'b011;
	13'd2319: q = 3'b011;
	13'd2320: q = 3'b011;
	13'd2321: q = 3'b011;
	13'd2322: q = 3'b011;
	13'd2323: q = 3'b011;
	13'd2324: q = 3'b011;
	13'd2325: q = 3'b011;
	13'd2326: q = 3'b011;
	13'd2327: q = 3'b011;
	13'd2328: q = 3'b011;
	13'd2329: q = 3'b011;
	13'd2330: q = 3'b011;
	13'd2331: q = 3'b011;
	13'd2332: q = 3'b011;
	13'd2333: q = 3'b011;
	13'd2334: q = 3'b000;
	13'd2335: q = 3'b000;
	13'd2336: q = 3'b111;
	13'd2337: q = 3'b111;
	13'd2338: q = 3'b011;
	13'd2339: q = 3'b011;
	13'd2340: q = 3'b011;
	13'd2341: q = 3'b011;
	13'd2342: q = 3'b011;
	13'd2343: q = 3'b011;
	13'd2344: q = 3'b011;
	13'd2345: q = 3'b011;
	13'd2346: q = 3'b011;
	13'd2347: q = 3'b011;
	13'd2348: q = 3'b011;
	13'd2349: q = 3'b011;
	13'd2350: q = 3'b011;
	13'd2351: q = 3'b011;
	13'd2352: q = 3'b011;
	13'd2353: q = 3'b011;
	13'd2354: q = 3'b011;
	13'd2355: q = 3'b011;
	13'd2356: q = 3'b011;
	13'd2357: q = 3'b011;
	13'd2358: q = 3'b011;
	13'd2359: q = 3'b011;
	13'd2360: q = 3'b011;
	13'd2361: q = 3'b011;
	13'd2362: q = 3'b011;
	13'd2363: q = 3'b011;
	13'd2364: q = 3'b011;
	13'd2365: q = 3'b011;
	13'd2366: q = 3'b000;
	13'd2367: q = 3'b000;
	13'd2368: q = 3'b000;
	13'd2369: q = 3'b000;
	13'd2370: q = 3'b000;
	13'd2371: q = 3'b000;
	13'd2372: q = 3'b000;
	13'd2373: q = 3'b000;
	13'd2374: q = 3'b000;
	13'd2375: q = 3'b000;
	13'd2376: q = 3'b000;
	13'd2377: q = 3'b000;
	13'd2378: q = 3'b000;
	13'd2379: q = 3'b000;
	13'd2380: q = 3'b000;
	13'd2381: q = 3'b000;
	13'd2382: q = 3'b000;
	13'd2383: q = 3'b000;
	13'd2384: q = 3'b000;
	13'd2385: q = 3'b000;
	13'd2386: q = 3'b000;
	13'd2387: q = 3'b000;
	13'd2388: q = 3'b000;
	13'd2389: q = 3'b000;
	13'd2390: q = 3'b000;
	13'd2391: q = 3'b000;
	13'd2392: q = 3'b000;
	13'd2393: q = 3'b000;
	13'd2394: q = 3'b000;
	13'd2395: q = 3'b000;
	13'd2396: q = 3'b000;
	13'd2397: q = 3'b000;
	13'd2398: q = 3'b000;
	13'd2399: q = 3'b000;
	13'd2400: q = 3'b000;
	13'd2401: q = 3'b000;
	13'd2402: q = 3'b000;
	13'd2403: q = 3'b000;
	13'd2404: q = 3'b000;
	13'd2405: q = 3'b000;
	13'd2406: q = 3'b000;
	13'd2407: q = 3'b000;
	13'd2408: q = 3'b000;
	13'd2409: q = 3'b000;
	13'd2410: q = 3'b000;
	13'd2411: q = 3'b000;
	13'd2412: q = 3'b000;
	13'd2413: q = 3'b000;
	13'd2414: q = 3'b000;
	13'd2415: q = 3'b000;
	13'd2416: q = 3'b000;
	13'd2417: q = 3'b000;
	13'd2418: q = 3'b000;
	13'd2419: q = 3'b000;
	13'd2420: q = 3'b000;
	13'd2421: q = 3'b000;
	13'd2422: q = 3'b000;
	13'd2423: q = 3'b000;
	13'd2424: q = 3'b000;
	13'd2425: q = 3'b000;
	13'd2426: q = 3'b000;
	13'd2427: q = 3'b000;
	13'd2428: q = 3'b000;
	13'd2429: q = 3'b000;
	13'd2430: q = 3'b000;
	13'd2431: q = 3'b000;
	13'd2432: q = 3'b111;
	13'd2433: q = 3'b111;
	13'd2434: q = 3'b111;
	13'd2435: q = 3'b111;
	13'd2436: q = 3'b111;
	13'd2437: q = 3'b111;
	13'd2438: q = 3'b111;
	13'd2439: q = 3'b111;
	13'd2440: q = 3'b111;
	13'd2441: q = 3'b111;
	13'd2442: q = 3'b000;
	13'd2443: q = 3'b000;
	13'd2444: q = 3'b000;
	13'd2445: q = 3'b000;
	13'd2446: q = 3'b111;
	13'd2447: q = 3'b111;
	13'd2448: q = 3'b111;
	13'd2449: q = 3'b111;
	13'd2450: q = 3'b111;
	13'd2451: q = 3'b111;
	13'd2452: q = 3'b111;
	13'd2453: q = 3'b111;
	13'd2454: q = 3'b111;
	13'd2455: q = 3'b111;
	13'd2456: q = 3'b111;
	13'd2457: q = 3'b111;
	13'd2458: q = 3'b111;
	13'd2459: q = 3'b111;
	13'd2460: q = 3'b111;
	13'd2461: q = 3'b111;
	13'd2462: q = 3'b111;
	13'd2463: q = 3'b111;
	13'd2464: q = 3'b111;
	13'd2465: q = 3'b111;
	13'd2466: q = 3'b111;
	13'd2467: q = 3'b111;
	13'd2468: q = 3'b111;
	13'd2469: q = 3'b111;
	13'd2470: q = 3'b111;
	13'd2471: q = 3'b111;
	13'd2472: q = 3'b111;
	13'd2473: q = 3'b111;
	13'd2474: q = 3'b000;
	13'd2475: q = 3'b000;
	13'd2476: q = 3'b000;
	13'd2477: q = 3'b000;
	13'd2478: q = 3'b111;
	13'd2479: q = 3'b111;
	13'd2480: q = 3'b111;
	13'd2481: q = 3'b111;
	13'd2482: q = 3'b111;
	13'd2483: q = 3'b111;
	13'd2484: q = 3'b111;
	13'd2485: q = 3'b111;
	13'd2486: q = 3'b111;
	13'd2487: q = 3'b111;
	13'd2488: q = 3'b111;
	13'd2489: q = 3'b111;
	13'd2490: q = 3'b111;
	13'd2491: q = 3'b111;
	13'd2492: q = 3'b111;
	13'd2493: q = 3'b111;
	13'd2494: q = 3'b111;
	13'd2495: q = 3'b111;
	13'd2496: q = 3'b011;
	13'd2497: q = 3'b011;
	13'd2498: q = 3'b011;
	13'd2499: q = 3'b011;
	13'd2500: q = 3'b011;
	13'd2501: q = 3'b011;
	13'd2502: q = 3'b011;
	13'd2503: q = 3'b011;
	13'd2504: q = 3'b011;
	13'd2505: q = 3'b011;
	13'd2506: q = 3'b000;
	13'd2507: q = 3'b000;
	13'd2508: q = 3'b111;
	13'd2509: q = 3'b111;
	13'd2510: q = 3'b011;
	13'd2511: q = 3'b011;
	13'd2512: q = 3'b011;
	13'd2513: q = 3'b011;
	13'd2514: q = 3'b011;
	13'd2515: q = 3'b011;
	13'd2516: q = 3'b011;
	13'd2517: q = 3'b011;
	13'd2518: q = 3'b011;
	13'd2519: q = 3'b011;
	13'd2520: q = 3'b011;
	13'd2521: q = 3'b011;
	13'd2522: q = 3'b011;
	13'd2523: q = 3'b011;
	13'd2524: q = 3'b011;
	13'd2525: q = 3'b011;
	13'd2526: q = 3'b011;
	13'd2527: q = 3'b011;
	13'd2528: q = 3'b011;
	13'd2529: q = 3'b011;
	13'd2530: q = 3'b011;
	13'd2531: q = 3'b011;
	13'd2532: q = 3'b011;
	13'd2533: q = 3'b011;
	13'd2534: q = 3'b011;
	13'd2535: q = 3'b011;
	13'd2536: q = 3'b011;
	13'd2537: q = 3'b011;
	13'd2538: q = 3'b000;
	13'd2539: q = 3'b000;
	13'd2540: q = 3'b111;
	13'd2541: q = 3'b111;
	13'd2542: q = 3'b011;
	13'd2543: q = 3'b011;
	13'd2544: q = 3'b011;
	13'd2545: q = 3'b011;
	13'd2546: q = 3'b011;
	13'd2547: q = 3'b011;
	13'd2548: q = 3'b011;
	13'd2549: q = 3'b011;
	13'd2550: q = 3'b011;
	13'd2551: q = 3'b011;
	13'd2552: q = 3'b011;
	13'd2553: q = 3'b011;
	13'd2554: q = 3'b011;
	13'd2555: q = 3'b011;
	13'd2556: q = 3'b011;
	13'd2557: q = 3'b011;
	13'd2558: q = 3'b011;
	13'd2559: q = 3'b011;
	13'd2560: q = 3'b011;
	13'd2561: q = 3'b011;
	13'd2562: q = 3'b011;
	13'd2563: q = 3'b011;
	13'd2564: q = 3'b011;
	13'd2565: q = 3'b011;
	13'd2566: q = 3'b011;
	13'd2567: q = 3'b011;
	13'd2568: q = 3'b011;
	13'd2569: q = 3'b011;
	13'd2570: q = 3'b000;
	13'd2571: q = 3'b000;
	13'd2572: q = 3'b111;
	13'd2573: q = 3'b111;
	13'd2574: q = 3'b011;
	13'd2575: q = 3'b011;
	13'd2576: q = 3'b011;
	13'd2577: q = 3'b011;
	13'd2578: q = 3'b011;
	13'd2579: q = 3'b011;
	13'd2580: q = 3'b011;
	13'd2581: q = 3'b011;
	13'd2582: q = 3'b011;
	13'd2583: q = 3'b011;
	13'd2584: q = 3'b011;
	13'd2585: q = 3'b011;
	13'd2586: q = 3'b011;
	13'd2587: q = 3'b011;
	13'd2588: q = 3'b011;
	13'd2589: q = 3'b011;
	13'd2590: q = 3'b011;
	13'd2591: q = 3'b011;
	13'd2592: q = 3'b011;
	13'd2593: q = 3'b011;
	13'd2594: q = 3'b011;
	13'd2595: q = 3'b011;
	13'd2596: q = 3'b011;
	13'd2597: q = 3'b011;
	13'd2598: q = 3'b011;
	13'd2599: q = 3'b011;
	13'd2600: q = 3'b011;
	13'd2601: q = 3'b011;
	13'd2602: q = 3'b000;
	13'd2603: q = 3'b000;
	13'd2604: q = 3'b111;
	13'd2605: q = 3'b111;
	13'd2606: q = 3'b011;
	13'd2607: q = 3'b011;
	13'd2608: q = 3'b011;
	13'd2609: q = 3'b011;
	13'd2610: q = 3'b011;
	13'd2611: q = 3'b011;
	13'd2612: q = 3'b011;
	13'd2613: q = 3'b011;
	13'd2614: q = 3'b011;
	13'd2615: q = 3'b011;
	13'd2616: q = 3'b011;
	13'd2617: q = 3'b011;
	13'd2618: q = 3'b011;
	13'd2619: q = 3'b011;
	13'd2620: q = 3'b011;
	13'd2621: q = 3'b011;
	13'd2622: q = 3'b011;
	13'd2623: q = 3'b011;
	13'd2624: q = 3'b011;
	13'd2625: q = 3'b011;
	13'd2626: q = 3'b011;
	13'd2627: q = 3'b011;
	13'd2628: q = 3'b011;
	13'd2629: q = 3'b011;
	13'd2630: q = 3'b011;
	13'd2631: q = 3'b011;
	13'd2632: q = 3'b011;
	13'd2633: q = 3'b011;
	13'd2634: q = 3'b000;
	13'd2635: q = 3'b000;
	13'd2636: q = 3'b111;
	13'd2637: q = 3'b111;
	13'd2638: q = 3'b011;
	13'd2639: q = 3'b011;
	13'd2640: q = 3'b011;
	13'd2641: q = 3'b011;
	13'd2642: q = 3'b011;
	13'd2643: q = 3'b011;
	13'd2644: q = 3'b011;
	13'd2645: q = 3'b011;
	13'd2646: q = 3'b011;
	13'd2647: q = 3'b011;
	13'd2648: q = 3'b011;
	13'd2649: q = 3'b011;
	13'd2650: q = 3'b011;
	13'd2651: q = 3'b011;
	13'd2652: q = 3'b011;
	13'd2653: q = 3'b011;
	13'd2654: q = 3'b011;
	13'd2655: q = 3'b011;
	13'd2656: q = 3'b011;
	13'd2657: q = 3'b011;
	13'd2658: q = 3'b011;
	13'd2659: q = 3'b011;
	13'd2660: q = 3'b011;
	13'd2661: q = 3'b011;
	13'd2662: q = 3'b011;
	13'd2663: q = 3'b011;
	13'd2664: q = 3'b011;
	13'd2665: q = 3'b011;
	13'd2666: q = 3'b000;
	13'd2667: q = 3'b000;
	13'd2668: q = 3'b111;
	13'd2669: q = 3'b111;
	13'd2670: q = 3'b011;
	13'd2671: q = 3'b011;
	13'd2672: q = 3'b011;
	13'd2673: q = 3'b011;
	13'd2674: q = 3'b011;
	13'd2675: q = 3'b011;
	13'd2676: q = 3'b011;
	13'd2677: q = 3'b011;
	13'd2678: q = 3'b011;
	13'd2679: q = 3'b011;
	13'd2680: q = 3'b011;
	13'd2681: q = 3'b011;
	13'd2682: q = 3'b011;
	13'd2683: q = 3'b011;
	13'd2684: q = 3'b011;
	13'd2685: q = 3'b011;
	13'd2686: q = 3'b011;
	13'd2687: q = 3'b011;
	13'd2688: q = 3'b000;
	13'd2689: q = 3'b000;
	13'd2690: q = 3'b000;
	13'd2691: q = 3'b000;
	13'd2692: q = 3'b000;
	13'd2693: q = 3'b000;
	13'd2694: q = 3'b000;
	13'd2695: q = 3'b000;
	13'd2696: q = 3'b000;
	13'd2697: q = 3'b000;
	13'd2698: q = 3'b000;
	13'd2699: q = 3'b000;
	13'd2700: q = 3'b000;
	13'd2701: q = 3'b000;
	13'd2702: q = 3'b000;
	13'd2703: q = 3'b000;
	13'd2704: q = 3'b000;
	13'd2705: q = 3'b000;
	13'd2706: q = 3'b000;
	13'd2707: q = 3'b000;
	13'd2708: q = 3'b000;
	13'd2709: q = 3'b000;
	13'd2710: q = 3'b000;
	13'd2711: q = 3'b000;
	13'd2712: q = 3'b000;
	13'd2713: q = 3'b000;
	13'd2714: q = 3'b000;
	13'd2715: q = 3'b000;
	13'd2716: q = 3'b000;
	13'd2717: q = 3'b000;
	13'd2718: q = 3'b000;
	13'd2719: q = 3'b000;
	13'd2720: q = 3'b000;
	13'd2721: q = 3'b000;
	13'd2722: q = 3'b000;
	13'd2723: q = 3'b000;
	13'd2724: q = 3'b000;
	13'd2725: q = 3'b000;
	13'd2726: q = 3'b000;
	13'd2727: q = 3'b000;
	13'd2728: q = 3'b000;
	13'd2729: q = 3'b000;
	13'd2730: q = 3'b000;
	13'd2731: q = 3'b000;
	13'd2732: q = 3'b000;
	13'd2733: q = 3'b000;
	13'd2734: q = 3'b000;
	13'd2735: q = 3'b000;
	13'd2736: q = 3'b000;
	13'd2737: q = 3'b000;
	13'd2738: q = 3'b000;
	13'd2739: q = 3'b000;
	13'd2740: q = 3'b000;
	13'd2741: q = 3'b000;
	13'd2742: q = 3'b000;
	13'd2743: q = 3'b000;
	13'd2744: q = 3'b000;
	13'd2745: q = 3'b000;
	13'd2746: q = 3'b000;
	13'd2747: q = 3'b000;
	13'd2748: q = 3'b000;
	13'd2749: q = 3'b000;
	13'd2750: q = 3'b000;
	13'd2751: q = 3'b000;
	13'd2752: q = 3'b111;
	13'd2753: q = 3'b111;
	13'd2754: q = 3'b111;
	13'd2755: q = 3'b111;
	13'd2756: q = 3'b111;
	13'd2757: q = 3'b111;
	13'd2758: q = 3'b111;
	13'd2759: q = 3'b111;
	13'd2760: q = 3'b111;
	13'd2761: q = 3'b111;
	13'd2762: q = 3'b111;
	13'd2763: q = 3'b111;
	13'd2764: q = 3'b111;
	13'd2765: q = 3'b111;
	13'd2766: q = 3'b111;
	13'd2767: q = 3'b111;
	13'd2768: q = 3'b111;
	13'd2769: q = 3'b111;
	13'd2770: q = 3'b000;
	13'd2771: q = 3'b000;
	13'd2772: q = 3'b000;
	13'd2773: q = 3'b000;
	13'd2774: q = 3'b111;
	13'd2775: q = 3'b111;
	13'd2776: q = 3'b111;
	13'd2777: q = 3'b111;
	13'd2778: q = 3'b111;
	13'd2779: q = 3'b111;
	13'd2780: q = 3'b111;
	13'd2781: q = 3'b111;
	13'd2782: q = 3'b111;
	13'd2783: q = 3'b111;
	13'd2784: q = 3'b111;
	13'd2785: q = 3'b111;
	13'd2786: q = 3'b111;
	13'd2787: q = 3'b111;
	13'd2788: q = 3'b111;
	13'd2789: q = 3'b111;
	13'd2790: q = 3'b111;
	13'd2791: q = 3'b111;
	13'd2792: q = 3'b111;
	13'd2793: q = 3'b111;
	13'd2794: q = 3'b111;
	13'd2795: q = 3'b111;
	13'd2796: q = 3'b111;
	13'd2797: q = 3'b111;
	13'd2798: q = 3'b111;
	13'd2799: q = 3'b111;
	13'd2800: q = 3'b111;
	13'd2801: q = 3'b111;
	13'd2802: q = 3'b000;
	13'd2803: q = 3'b000;
	13'd2804: q = 3'b000;
	13'd2805: q = 3'b000;
	13'd2806: q = 3'b111;
	13'd2807: q = 3'b111;
	13'd2808: q = 3'b111;
	13'd2809: q = 3'b111;
	13'd2810: q = 3'b111;
	13'd2811: q = 3'b111;
	13'd2812: q = 3'b111;
	13'd2813: q = 3'b111;
	13'd2814: q = 3'b111;
	13'd2815: q = 3'b111;
	13'd2816: q = 3'b011;
	13'd2817: q = 3'b011;
	13'd2818: q = 3'b011;
	13'd2819: q = 3'b011;
	13'd2820: q = 3'b011;
	13'd2821: q = 3'b011;
	13'd2822: q = 3'b011;
	13'd2823: q = 3'b011;
	13'd2824: q = 3'b011;
	13'd2825: q = 3'b011;
	13'd2826: q = 3'b011;
	13'd2827: q = 3'b011;
	13'd2828: q = 3'b011;
	13'd2829: q = 3'b011;
	13'd2830: q = 3'b011;
	13'd2831: q = 3'b011;
	13'd2832: q = 3'b011;
	13'd2833: q = 3'b011;
	13'd2834: q = 3'b000;
	13'd2835: q = 3'b000;
	13'd2836: q = 3'b111;
	13'd2837: q = 3'b111;
	13'd2838: q = 3'b011;
	13'd2839: q = 3'b011;
	13'd2840: q = 3'b011;
	13'd2841: q = 3'b011;
	13'd2842: q = 3'b011;
	13'd2843: q = 3'b011;
	13'd2844: q = 3'b011;
	13'd2845: q = 3'b011;
	13'd2846: q = 3'b011;
	13'd2847: q = 3'b011;
	13'd2848: q = 3'b011;
	13'd2849: q = 3'b011;
	13'd2850: q = 3'b011;
	13'd2851: q = 3'b011;
	13'd2852: q = 3'b011;
	13'd2853: q = 3'b011;
	13'd2854: q = 3'b011;
	13'd2855: q = 3'b011;
	13'd2856: q = 3'b011;
	13'd2857: q = 3'b011;
	13'd2858: q = 3'b011;
	13'd2859: q = 3'b011;
	13'd2860: q = 3'b011;
	13'd2861: q = 3'b011;
	13'd2862: q = 3'b011;
	13'd2863: q = 3'b011;
	13'd2864: q = 3'b011;
	13'd2865: q = 3'b011;
	13'd2866: q = 3'b000;
	13'd2867: q = 3'b000;
	13'd2868: q = 3'b111;
	13'd2869: q = 3'b111;
	13'd2870: q = 3'b011;
	13'd2871: q = 3'b011;
	13'd2872: q = 3'b011;
	13'd2873: q = 3'b011;
	13'd2874: q = 3'b011;
	13'd2875: q = 3'b011;
	13'd2876: q = 3'b011;
	13'd2877: q = 3'b011;
	13'd2878: q = 3'b011;
	13'd2879: q = 3'b011;
	13'd2880: q = 3'b011;
	13'd2881: q = 3'b011;
	13'd2882: q = 3'b011;
	13'd2883: q = 3'b011;
	13'd2884: q = 3'b011;
	13'd2885: q = 3'b011;
	13'd2886: q = 3'b011;
	13'd2887: q = 3'b011;
	13'd2888: q = 3'b011;
	13'd2889: q = 3'b011;
	13'd2890: q = 3'b011;
	13'd2891: q = 3'b011;
	13'd2892: q = 3'b011;
	13'd2893: q = 3'b011;
	13'd2894: q = 3'b011;
	13'd2895: q = 3'b011;
	13'd2896: q = 3'b011;
	13'd2897: q = 3'b011;
	13'd2898: q = 3'b000;
	13'd2899: q = 3'b000;
	13'd2900: q = 3'b111;
	13'd2901: q = 3'b111;
	13'd2902: q = 3'b011;
	13'd2903: q = 3'b011;
	13'd2904: q = 3'b011;
	13'd2905: q = 3'b011;
	13'd2906: q = 3'b011;
	13'd2907: q = 3'b011;
	13'd2908: q = 3'b011;
	13'd2909: q = 3'b011;
	13'd2910: q = 3'b011;
	13'd2911: q = 3'b011;
	13'd2912: q = 3'b011;
	13'd2913: q = 3'b011;
	13'd2914: q = 3'b011;
	13'd2915: q = 3'b011;
	13'd2916: q = 3'b011;
	13'd2917: q = 3'b011;
	13'd2918: q = 3'b011;
	13'd2919: q = 3'b011;
	13'd2920: q = 3'b011;
	13'd2921: q = 3'b011;
	13'd2922: q = 3'b011;
	13'd2923: q = 3'b011;
	13'd2924: q = 3'b011;
	13'd2925: q = 3'b011;
	13'd2926: q = 3'b011;
	13'd2927: q = 3'b011;
	13'd2928: q = 3'b011;
	13'd2929: q = 3'b011;
	13'd2930: q = 3'b000;
	13'd2931: q = 3'b000;
	13'd2932: q = 3'b111;
	13'd2933: q = 3'b111;
	13'd2934: q = 3'b011;
	13'd2935: q = 3'b011;
	13'd2936: q = 3'b011;
	13'd2937: q = 3'b011;
	13'd2938: q = 3'b011;
	13'd2939: q = 3'b011;
	13'd2940: q = 3'b011;
	13'd2941: q = 3'b011;
	13'd2942: q = 3'b011;
	13'd2943: q = 3'b011;
	13'd2944: q = 3'b011;
	13'd2945: q = 3'b011;
	13'd2946: q = 3'b011;
	13'd2947: q = 3'b011;
	13'd2948: q = 3'b011;
	13'd2949: q = 3'b011;
	13'd2950: q = 3'b011;
	13'd2951: q = 3'b011;
	13'd2952: q = 3'b011;
	13'd2953: q = 3'b011;
	13'd2954: q = 3'b011;
	13'd2955: q = 3'b011;
	13'd2956: q = 3'b011;
	13'd2957: q = 3'b011;
	13'd2958: q = 3'b011;
	13'd2959: q = 3'b011;
	13'd2960: q = 3'b011;
	13'd2961: q = 3'b011;
	13'd2962: q = 3'b000;
	13'd2963: q = 3'b000;
	13'd2964: q = 3'b111;
	13'd2965: q = 3'b111;
	13'd2966: q = 3'b011;
	13'd2967: q = 3'b011;
	13'd2968: q = 3'b011;
	13'd2969: q = 3'b011;
	13'd2970: q = 3'b011;
	13'd2971: q = 3'b011;
	13'd2972: q = 3'b011;
	13'd2973: q = 3'b011;
	13'd2974: q = 3'b011;
	13'd2975: q = 3'b011;
	13'd2976: q = 3'b011;
	13'd2977: q = 3'b011;
	13'd2978: q = 3'b011;
	13'd2979: q = 3'b011;
	13'd2980: q = 3'b011;
	13'd2981: q = 3'b011;
	13'd2982: q = 3'b011;
	13'd2983: q = 3'b011;
	13'd2984: q = 3'b011;
	13'd2985: q = 3'b011;
	13'd2986: q = 3'b011;
	13'd2987: q = 3'b011;
	13'd2988: q = 3'b011;
	13'd2989: q = 3'b011;
	13'd2990: q = 3'b011;
	13'd2991: q = 3'b011;
	13'd2992: q = 3'b011;
	13'd2993: q = 3'b011;
	13'd2994: q = 3'b000;
	13'd2995: q = 3'b000;
	13'd2996: q = 3'b111;
	13'd2997: q = 3'b111;
	13'd2998: q = 3'b011;
	13'd2999: q = 3'b011;
	13'd3000: q = 3'b011;
	13'd3001: q = 3'b011;
	13'd3002: q = 3'b011;
	13'd3003: q = 3'b011;
	13'd3004: q = 3'b011;
	13'd3005: q = 3'b011;
	13'd3006: q = 3'b011;
	13'd3007: q = 3'b011;
	13'd3008: q = 3'b000;
	13'd3009: q = 3'b000;
	13'd3010: q = 3'b000;
	13'd3011: q = 3'b000;
	13'd3012: q = 3'b000;
	13'd3013: q = 3'b000;
	13'd3014: q = 3'b000;
	13'd3015: q = 3'b000;
	13'd3016: q = 3'b000;
	13'd3017: q = 3'b000;
	13'd3018: q = 3'b000;
	13'd3019: q = 3'b000;
	13'd3020: q = 3'b000;
	13'd3021: q = 3'b000;
	13'd3022: q = 3'b000;
	13'd3023: q = 3'b000;
	13'd3024: q = 3'b000;
	13'd3025: q = 3'b000;
	13'd3026: q = 3'b000;
	13'd3027: q = 3'b000;
	13'd3028: q = 3'b000;
	13'd3029: q = 3'b000;
	13'd3030: q = 3'b000;
	13'd3031: q = 3'b000;
	13'd3032: q = 3'b000;
	13'd3033: q = 3'b000;
	13'd3034: q = 3'b000;
	13'd3035: q = 3'b000;
	13'd3036: q = 3'b000;
	13'd3037: q = 3'b000;
	13'd3038: q = 3'b000;
	13'd3039: q = 3'b000;
	13'd3040: q = 3'b000;
	13'd3041: q = 3'b000;
	13'd3042: q = 3'b000;
	13'd3043: q = 3'b000;
	13'd3044: q = 3'b000;
	13'd3045: q = 3'b000;
	13'd3046: q = 3'b000;
	13'd3047: q = 3'b000;
	13'd3048: q = 3'b000;
	13'd3049: q = 3'b000;
	13'd3050: q = 3'b000;
	13'd3051: q = 3'b000;
	13'd3052: q = 3'b000;
	13'd3053: q = 3'b000;
	13'd3054: q = 3'b000;
	13'd3055: q = 3'b000;
	13'd3056: q = 3'b000;
	13'd3057: q = 3'b000;
	13'd3058: q = 3'b000;
	13'd3059: q = 3'b000;
	13'd3060: q = 3'b000;
	13'd3061: q = 3'b000;
	13'd3062: q = 3'b000;
	13'd3063: q = 3'b000;
	13'd3064: q = 3'b000;
	13'd3065: q = 3'b000;
	13'd3066: q = 3'b000;
	13'd3067: q = 3'b000;
	13'd3068: q = 3'b000;
	13'd3069: q = 3'b000;
	13'd3070: q = 3'b000;
	13'd3071: q = 3'b000;
	13'd3072: q = 3'b011;
	13'd3073: q = 3'b011;
	13'd3074: q = 3'b111;
	13'd3075: q = 3'b111;
	13'd3076: q = 3'b111;
	13'd3077: q = 3'b111;
	13'd3078: q = 3'b111;
	13'd3079: q = 3'b111;
	13'd3080: q = 3'b111;
	13'd3081: q = 3'b111;
	13'd3082: q = 3'b111;
	13'd3083: q = 3'b111;
	13'd3084: q = 3'b111;
	13'd3085: q = 3'b111;
	13'd3086: q = 3'b111;
	13'd3087: q = 3'b111;
	13'd3088: q = 3'b111;
	13'd3089: q = 3'b111;
	13'd3090: q = 3'b111;
	13'd3091: q = 3'b111;
	13'd3092: q = 3'b111;
	13'd3093: q = 3'b111;
	13'd3094: q = 3'b111;
	13'd3095: q = 3'b111;
	13'd3096: q = 3'b111;
	13'd3097: q = 3'b111;
	13'd3098: q = 3'b111;
	13'd3099: q = 3'b111;
	13'd3100: q = 3'b111;
	13'd3101: q = 3'b111;
	13'd3102: q = 3'b000;
	13'd3103: q = 3'b000;
	13'd3104: q = 3'b011;
	13'd3105: q = 3'b011;
	13'd3106: q = 3'b111;
	13'd3107: q = 3'b111;
	13'd3108: q = 3'b111;
	13'd3109: q = 3'b111;
	13'd3110: q = 3'b111;
	13'd3111: q = 3'b111;
	13'd3112: q = 3'b111;
	13'd3113: q = 3'b111;
	13'd3114: q = 3'b111;
	13'd3115: q = 3'b111;
	13'd3116: q = 3'b111;
	13'd3117: q = 3'b111;
	13'd3118: q = 3'b111;
	13'd3119: q = 3'b111;
	13'd3120: q = 3'b111;
	13'd3121: q = 3'b111;
	13'd3122: q = 3'b111;
	13'd3123: q = 3'b111;
	13'd3124: q = 3'b111;
	13'd3125: q = 3'b111;
	13'd3126: q = 3'b111;
	13'd3127: q = 3'b111;
	13'd3128: q = 3'b111;
	13'd3129: q = 3'b111;
	13'd3130: q = 3'b111;
	13'd3131: q = 3'b111;
	13'd3132: q = 3'b111;
	13'd3133: q = 3'b111;
	13'd3134: q = 3'b000;
	13'd3135: q = 3'b000;
	13'd3136: q = 3'b111;
	13'd3137: q = 3'b111;
	13'd3138: q = 3'b100;
	13'd3139: q = 3'b100;
	13'd3140: q = 3'b100;
	13'd3141: q = 3'b100;
	13'd3142: q = 3'b100;
	13'd3143: q = 3'b100;
	13'd3144: q = 3'b100;
	13'd3145: q = 3'b100;
	13'd3146: q = 3'b100;
	13'd3147: q = 3'b100;
	13'd3148: q = 3'b100;
	13'd3149: q = 3'b100;
	13'd3150: q = 3'b100;
	13'd3151: q = 3'b100;
	13'd3152: q = 3'b100;
	13'd3153: q = 3'b100;
	13'd3154: q = 3'b100;
	13'd3155: q = 3'b100;
	13'd3156: q = 3'b100;
	13'd3157: q = 3'b100;
	13'd3158: q = 3'b100;
	13'd3159: q = 3'b100;
	13'd3160: q = 3'b100;
	13'd3161: q = 3'b100;
	13'd3162: q = 3'b100;
	13'd3163: q = 3'b100;
	13'd3164: q = 3'b100;
	13'd3165: q = 3'b100;
	13'd3166: q = 3'b000;
	13'd3167: q = 3'b000;
	13'd3168: q = 3'b111;
	13'd3169: q = 3'b111;
	13'd3170: q = 3'b100;
	13'd3171: q = 3'b100;
	13'd3172: q = 3'b100;
	13'd3173: q = 3'b100;
	13'd3174: q = 3'b100;
	13'd3175: q = 3'b100;
	13'd3176: q = 3'b100;
	13'd3177: q = 3'b100;
	13'd3178: q = 3'b100;
	13'd3179: q = 3'b100;
	13'd3180: q = 3'b100;
	13'd3181: q = 3'b100;
	13'd3182: q = 3'b100;
	13'd3183: q = 3'b100;
	13'd3184: q = 3'b100;
	13'd3185: q = 3'b100;
	13'd3186: q = 3'b100;
	13'd3187: q = 3'b100;
	13'd3188: q = 3'b100;
	13'd3189: q = 3'b100;
	13'd3190: q = 3'b100;
	13'd3191: q = 3'b100;
	13'd3192: q = 3'b100;
	13'd3193: q = 3'b100;
	13'd3194: q = 3'b100;
	13'd3195: q = 3'b100;
	13'd3196: q = 3'b100;
	13'd3197: q = 3'b100;
	13'd3198: q = 3'b000;
	13'd3199: q = 3'b000;
	13'd3200: q = 3'b111;
	13'd3201: q = 3'b111;
	13'd3202: q = 3'b100;
	13'd3203: q = 3'b100;
	13'd3204: q = 3'b100;
	13'd3205: q = 3'b100;
	13'd3206: q = 3'b100;
	13'd3207: q = 3'b100;
	13'd3208: q = 3'b100;
	13'd3209: q = 3'b100;
	13'd3210: q = 3'b100;
	13'd3211: q = 3'b100;
	13'd3212: q = 3'b100;
	13'd3213: q = 3'b100;
	13'd3214: q = 3'b100;
	13'd3215: q = 3'b100;
	13'd3216: q = 3'b100;
	13'd3217: q = 3'b100;
	13'd3218: q = 3'b100;
	13'd3219: q = 3'b100;
	13'd3220: q = 3'b100;
	13'd3221: q = 3'b100;
	13'd3222: q = 3'b100;
	13'd3223: q = 3'b100;
	13'd3224: q = 3'b100;
	13'd3225: q = 3'b100;
	13'd3226: q = 3'b100;
	13'd3227: q = 3'b100;
	13'd3228: q = 3'b100;
	13'd3229: q = 3'b100;
	13'd3230: q = 3'b000;
	13'd3231: q = 3'b000;
	13'd3232: q = 3'b111;
	13'd3233: q = 3'b111;
	13'd3234: q = 3'b100;
	13'd3235: q = 3'b100;
	13'd3236: q = 3'b100;
	13'd3237: q = 3'b100;
	13'd3238: q = 3'b100;
	13'd3239: q = 3'b100;
	13'd3240: q = 3'b100;
	13'd3241: q = 3'b100;
	13'd3242: q = 3'b100;
	13'd3243: q = 3'b100;
	13'd3244: q = 3'b100;
	13'd3245: q = 3'b100;
	13'd3246: q = 3'b100;
	13'd3247: q = 3'b100;
	13'd3248: q = 3'b100;
	13'd3249: q = 3'b100;
	13'd3250: q = 3'b100;
	13'd3251: q = 3'b100;
	13'd3252: q = 3'b100;
	13'd3253: q = 3'b100;
	13'd3254: q = 3'b100;
	13'd3255: q = 3'b100;
	13'd3256: q = 3'b100;
	13'd3257: q = 3'b100;
	13'd3258: q = 3'b100;
	13'd3259: q = 3'b100;
	13'd3260: q = 3'b100;
	13'd3261: q = 3'b100;
	13'd3262: q = 3'b000;
	13'd3263: q = 3'b000;
	13'd3264: q = 3'b111;
	13'd3265: q = 3'b111;
	13'd3266: q = 3'b100;
	13'd3267: q = 3'b100;
	13'd3268: q = 3'b100;
	13'd3269: q = 3'b100;
	13'd3270: q = 3'b100;
	13'd3271: q = 3'b100;
	13'd3272: q = 3'b100;
	13'd3273: q = 3'b100;
	13'd3274: q = 3'b100;
	13'd3275: q = 3'b100;
	13'd3276: q = 3'b100;
	13'd3277: q = 3'b100;
	13'd3278: q = 3'b100;
	13'd3279: q = 3'b100;
	13'd3280: q = 3'b100;
	13'd3281: q = 3'b100;
	13'd3282: q = 3'b100;
	13'd3283: q = 3'b100;
	13'd3284: q = 3'b100;
	13'd3285: q = 3'b100;
	13'd3286: q = 3'b100;
	13'd3287: q = 3'b100;
	13'd3288: q = 3'b100;
	13'd3289: q = 3'b100;
	13'd3290: q = 3'b100;
	13'd3291: q = 3'b100;
	13'd3292: q = 3'b100;
	13'd3293: q = 3'b100;
	13'd3294: q = 3'b000;
	13'd3295: q = 3'b000;
	13'd3296: q = 3'b111;
	13'd3297: q = 3'b111;
	13'd3298: q = 3'b100;
	13'd3299: q = 3'b100;
	13'd3300: q = 3'b100;
	13'd3301: q = 3'b100;
	13'd3302: q = 3'b100;
	13'd3303: q = 3'b100;
	13'd3304: q = 3'b100;
	13'd3305: q = 3'b100;
	13'd3306: q = 3'b100;
	13'd3307: q = 3'b100;
	13'd3308: q = 3'b100;
	13'd3309: q = 3'b100;
	13'd3310: q = 3'b100;
	13'd3311: q = 3'b100;
	13'd3312: q = 3'b100;
	13'd3313: q = 3'b100;
	13'd3314: q = 3'b100;
	13'd3315: q = 3'b100;
	13'd3316: q = 3'b100;
	13'd3317: q = 3'b100;
	13'd3318: q = 3'b100;
	13'd3319: q = 3'b100;
	13'd3320: q = 3'b100;
	13'd3321: q = 3'b100;
	13'd3322: q = 3'b100;
	13'd3323: q = 3'b100;
	13'd3324: q = 3'b100;
	13'd3325: q = 3'b100;
	13'd3326: q = 3'b000;
	13'd3327: q = 3'b000;
	13'd3328: q = 3'b111;
	13'd3329: q = 3'b111;
	13'd3330: q = 3'b100;
	13'd3331: q = 3'b100;
	13'd3332: q = 3'b100;
	13'd3333: q = 3'b100;
	13'd3334: q = 3'b100;
	13'd3335: q = 3'b100;
	13'd3336: q = 3'b100;
	13'd3337: q = 3'b100;
	13'd3338: q = 3'b100;
	13'd3339: q = 3'b100;
	13'd3340: q = 3'b100;
	13'd3341: q = 3'b100;
	13'd3342: q = 3'b100;
	13'd3343: q = 3'b100;
	13'd3344: q = 3'b100;
	13'd3345: q = 3'b100;
	13'd3346: q = 3'b100;
	13'd3347: q = 3'b100;
	13'd3348: q = 3'b100;
	13'd3349: q = 3'b100;
	13'd3350: q = 3'b100;
	13'd3351: q = 3'b100;
	13'd3352: q = 3'b100;
	13'd3353: q = 3'b100;
	13'd3354: q = 3'b100;
	13'd3355: q = 3'b100;
	13'd3356: q = 3'b100;
	13'd3357: q = 3'b100;
	13'd3358: q = 3'b000;
	13'd3359: q = 3'b000;
	13'd3360: q = 3'b111;
	13'd3361: q = 3'b111;
	13'd3362: q = 3'b100;
	13'd3363: q = 3'b100;
	13'd3364: q = 3'b100;
	13'd3365: q = 3'b100;
	13'd3366: q = 3'b100;
	13'd3367: q = 3'b100;
	13'd3368: q = 3'b100;
	13'd3369: q = 3'b100;
	13'd3370: q = 3'b100;
	13'd3371: q = 3'b100;
	13'd3372: q = 3'b100;
	13'd3373: q = 3'b100;
	13'd3374: q = 3'b100;
	13'd3375: q = 3'b100;
	13'd3376: q = 3'b100;
	13'd3377: q = 3'b100;
	13'd3378: q = 3'b100;
	13'd3379: q = 3'b100;
	13'd3380: q = 3'b100;
	13'd3381: q = 3'b100;
	13'd3382: q = 3'b100;
	13'd3383: q = 3'b100;
	13'd3384: q = 3'b100;
	13'd3385: q = 3'b100;
	13'd3386: q = 3'b100;
	13'd3387: q = 3'b100;
	13'd3388: q = 3'b100;
	13'd3389: q = 3'b100;
	13'd3390: q = 3'b000;
	13'd3391: q = 3'b000;
	13'd3392: q = 3'b111;
	13'd3393: q = 3'b111;
	13'd3394: q = 3'b100;
	13'd3395: q = 3'b100;
	13'd3396: q = 3'b100;
	13'd3397: q = 3'b100;
	13'd3398: q = 3'b100;
	13'd3399: q = 3'b100;
	13'd3400: q = 3'b100;
	13'd3401: q = 3'b100;
	13'd3402: q = 3'b100;
	13'd3403: q = 3'b100;
	13'd3404: q = 3'b100;
	13'd3405: q = 3'b100;
	13'd3406: q = 3'b100;
	13'd3407: q = 3'b100;
	13'd3408: q = 3'b100;
	13'd3409: q = 3'b100;
	13'd3410: q = 3'b100;
	13'd3411: q = 3'b100;
	13'd3412: q = 3'b100;
	13'd3413: q = 3'b100;
	13'd3414: q = 3'b100;
	13'd3415: q = 3'b100;
	13'd3416: q = 3'b100;
	13'd3417: q = 3'b100;
	13'd3418: q = 3'b100;
	13'd3419: q = 3'b100;
	13'd3420: q = 3'b100;
	13'd3421: q = 3'b100;
	13'd3422: q = 3'b000;
	13'd3423: q = 3'b000;
	13'd3424: q = 3'b111;
	13'd3425: q = 3'b111;
	13'd3426: q = 3'b100;
	13'd3427: q = 3'b100;
	13'd3428: q = 3'b100;
	13'd3429: q = 3'b100;
	13'd3430: q = 3'b100;
	13'd3431: q = 3'b100;
	13'd3432: q = 3'b100;
	13'd3433: q = 3'b100;
	13'd3434: q = 3'b100;
	13'd3435: q = 3'b100;
	13'd3436: q = 3'b100;
	13'd3437: q = 3'b100;
	13'd3438: q = 3'b100;
	13'd3439: q = 3'b100;
	13'd3440: q = 3'b100;
	13'd3441: q = 3'b100;
	13'd3442: q = 3'b100;
	13'd3443: q = 3'b100;
	13'd3444: q = 3'b100;
	13'd3445: q = 3'b100;
	13'd3446: q = 3'b100;
	13'd3447: q = 3'b100;
	13'd3448: q = 3'b100;
	13'd3449: q = 3'b100;
	13'd3450: q = 3'b100;
	13'd3451: q = 3'b100;
	13'd3452: q = 3'b100;
	13'd3453: q = 3'b100;
	13'd3454: q = 3'b000;
	13'd3455: q = 3'b000;
	13'd3456: q = 3'b111;
	13'd3457: q = 3'b111;
	13'd3458: q = 3'b100;
	13'd3459: q = 3'b100;
	13'd3460: q = 3'b100;
	13'd3461: q = 3'b100;
	13'd3462: q = 3'b100;
	13'd3463: q = 3'b100;
	13'd3464: q = 3'b100;
	13'd3465: q = 3'b100;
	13'd3466: q = 3'b100;
	13'd3467: q = 3'b100;
	13'd3468: q = 3'b100;
	13'd3469: q = 3'b100;
	13'd3470: q = 3'b100;
	13'd3471: q = 3'b100;
	13'd3472: q = 3'b100;
	13'd3473: q = 3'b100;
	13'd3474: q = 3'b100;
	13'd3475: q = 3'b100;
	13'd3476: q = 3'b100;
	13'd3477: q = 3'b100;
	13'd3478: q = 3'b100;
	13'd3479: q = 3'b100;
	13'd3480: q = 3'b100;
	13'd3481: q = 3'b100;
	13'd3482: q = 3'b100;
	13'd3483: q = 3'b100;
	13'd3484: q = 3'b100;
	13'd3485: q = 3'b100;
	13'd3486: q = 3'b000;
	13'd3487: q = 3'b000;
	13'd3488: q = 3'b111;
	13'd3489: q = 3'b111;
	13'd3490: q = 3'b100;
	13'd3491: q = 3'b100;
	13'd3492: q = 3'b100;
	13'd3493: q = 3'b100;
	13'd3494: q = 3'b100;
	13'd3495: q = 3'b100;
	13'd3496: q = 3'b100;
	13'd3497: q = 3'b100;
	13'd3498: q = 3'b100;
	13'd3499: q = 3'b100;
	13'd3500: q = 3'b100;
	13'd3501: q = 3'b100;
	13'd3502: q = 3'b100;
	13'd3503: q = 3'b100;
	13'd3504: q = 3'b100;
	13'd3505: q = 3'b100;
	13'd3506: q = 3'b100;
	13'd3507: q = 3'b100;
	13'd3508: q = 3'b100;
	13'd3509: q = 3'b100;
	13'd3510: q = 3'b100;
	13'd3511: q = 3'b100;
	13'd3512: q = 3'b100;
	13'd3513: q = 3'b100;
	13'd3514: q = 3'b100;
	13'd3515: q = 3'b100;
	13'd3516: q = 3'b100;
	13'd3517: q = 3'b100;
	13'd3518: q = 3'b000;
	13'd3519: q = 3'b000;
	13'd3520: q = 3'b111;
	13'd3521: q = 3'b111;
	13'd3522: q = 3'b100;
	13'd3523: q = 3'b100;
	13'd3524: q = 3'b100;
	13'd3525: q = 3'b100;
	13'd3526: q = 3'b100;
	13'd3527: q = 3'b100;
	13'd3528: q = 3'b100;
	13'd3529: q = 3'b100;
	13'd3530: q = 3'b100;
	13'd3531: q = 3'b100;
	13'd3532: q = 3'b100;
	13'd3533: q = 3'b100;
	13'd3534: q = 3'b100;
	13'd3535: q = 3'b100;
	13'd3536: q = 3'b100;
	13'd3537: q = 3'b100;
	13'd3538: q = 3'b100;
	13'd3539: q = 3'b100;
	13'd3540: q = 3'b100;
	13'd3541: q = 3'b100;
	13'd3542: q = 3'b100;
	13'd3543: q = 3'b100;
	13'd3544: q = 3'b100;
	13'd3545: q = 3'b100;
	13'd3546: q = 3'b100;
	13'd3547: q = 3'b100;
	13'd3548: q = 3'b100;
	13'd3549: q = 3'b100;
	13'd3550: q = 3'b000;
	13'd3551: q = 3'b000;
	13'd3552: q = 3'b111;
	13'd3553: q = 3'b111;
	13'd3554: q = 3'b100;
	13'd3555: q = 3'b100;
	13'd3556: q = 3'b100;
	13'd3557: q = 3'b100;
	13'd3558: q = 3'b100;
	13'd3559: q = 3'b100;
	13'd3560: q = 3'b100;
	13'd3561: q = 3'b100;
	13'd3562: q = 3'b100;
	13'd3563: q = 3'b100;
	13'd3564: q = 3'b100;
	13'd3565: q = 3'b100;
	13'd3566: q = 3'b100;
	13'd3567: q = 3'b100;
	13'd3568: q = 3'b100;
	13'd3569: q = 3'b100;
	13'd3570: q = 3'b100;
	13'd3571: q = 3'b100;
	13'd3572: q = 3'b100;
	13'd3573: q = 3'b100;
	13'd3574: q = 3'b100;
	13'd3575: q = 3'b100;
	13'd3576: q = 3'b100;
	13'd3577: q = 3'b100;
	13'd3578: q = 3'b100;
	13'd3579: q = 3'b100;
	13'd3580: q = 3'b100;
	13'd3581: q = 3'b100;
	13'd3582: q = 3'b000;
	13'd3583: q = 3'b000;
	13'd3584: q = 3'b111;
	13'd3585: q = 3'b111;
	13'd3586: q = 3'b100;
	13'd3587: q = 3'b100;
	13'd3588: q = 3'b100;
	13'd3589: q = 3'b100;
	13'd3590: q = 3'b100;
	13'd3591: q = 3'b100;
	13'd3592: q = 3'b100;
	13'd3593: q = 3'b100;
	13'd3594: q = 3'b100;
	13'd3595: q = 3'b100;
	13'd3596: q = 3'b100;
	13'd3597: q = 3'b100;
	13'd3598: q = 3'b100;
	13'd3599: q = 3'b100;
	13'd3600: q = 3'b100;
	13'd3601: q = 3'b100;
	13'd3602: q = 3'b100;
	13'd3603: q = 3'b100;
	13'd3604: q = 3'b100;
	13'd3605: q = 3'b100;
	13'd3606: q = 3'b100;
	13'd3607: q = 3'b100;
	13'd3608: q = 3'b100;
	13'd3609: q = 3'b100;
	13'd3610: q = 3'b100;
	13'd3611: q = 3'b100;
	13'd3612: q = 3'b100;
	13'd3613: q = 3'b100;
	13'd3614: q = 3'b000;
	13'd3615: q = 3'b000;
	13'd3616: q = 3'b111;
	13'd3617: q = 3'b111;
	13'd3618: q = 3'b100;
	13'd3619: q = 3'b100;
	13'd3620: q = 3'b100;
	13'd3621: q = 3'b100;
	13'd3622: q = 3'b100;
	13'd3623: q = 3'b100;
	13'd3624: q = 3'b100;
	13'd3625: q = 3'b100;
	13'd3626: q = 3'b100;
	13'd3627: q = 3'b100;
	13'd3628: q = 3'b100;
	13'd3629: q = 3'b100;
	13'd3630: q = 3'b100;
	13'd3631: q = 3'b100;
	13'd3632: q = 3'b100;
	13'd3633: q = 3'b100;
	13'd3634: q = 3'b100;
	13'd3635: q = 3'b100;
	13'd3636: q = 3'b100;
	13'd3637: q = 3'b100;
	13'd3638: q = 3'b100;
	13'd3639: q = 3'b100;
	13'd3640: q = 3'b100;
	13'd3641: q = 3'b100;
	13'd3642: q = 3'b100;
	13'd3643: q = 3'b100;
	13'd3644: q = 3'b100;
	13'd3645: q = 3'b100;
	13'd3646: q = 3'b000;
	13'd3647: q = 3'b000;
	13'd3648: q = 3'b111;
	13'd3649: q = 3'b111;
	13'd3650: q = 3'b100;
	13'd3651: q = 3'b100;
	13'd3652: q = 3'b100;
	13'd3653: q = 3'b100;
	13'd3654: q = 3'b100;
	13'd3655: q = 3'b100;
	13'd3656: q = 3'b100;
	13'd3657: q = 3'b100;
	13'd3658: q = 3'b100;
	13'd3659: q = 3'b100;
	13'd3660: q = 3'b100;
	13'd3661: q = 3'b100;
	13'd3662: q = 3'b100;
	13'd3663: q = 3'b100;
	13'd3664: q = 3'b100;
	13'd3665: q = 3'b100;
	13'd3666: q = 3'b100;
	13'd3667: q = 3'b100;
	13'd3668: q = 3'b100;
	13'd3669: q = 3'b100;
	13'd3670: q = 3'b100;
	13'd3671: q = 3'b100;
	13'd3672: q = 3'b100;
	13'd3673: q = 3'b100;
	13'd3674: q = 3'b100;
	13'd3675: q = 3'b100;
	13'd3676: q = 3'b100;
	13'd3677: q = 3'b100;
	13'd3678: q = 3'b000;
	13'd3679: q = 3'b000;
	13'd3680: q = 3'b111;
	13'd3681: q = 3'b111;
	13'd3682: q = 3'b100;
	13'd3683: q = 3'b100;
	13'd3684: q = 3'b100;
	13'd3685: q = 3'b100;
	13'd3686: q = 3'b100;
	13'd3687: q = 3'b100;
	13'd3688: q = 3'b100;
	13'd3689: q = 3'b100;
	13'd3690: q = 3'b100;
	13'd3691: q = 3'b100;
	13'd3692: q = 3'b100;
	13'd3693: q = 3'b100;
	13'd3694: q = 3'b100;
	13'd3695: q = 3'b100;
	13'd3696: q = 3'b100;
	13'd3697: q = 3'b100;
	13'd3698: q = 3'b100;
	13'd3699: q = 3'b100;
	13'd3700: q = 3'b100;
	13'd3701: q = 3'b100;
	13'd3702: q = 3'b100;
	13'd3703: q = 3'b100;
	13'd3704: q = 3'b100;
	13'd3705: q = 3'b100;
	13'd3706: q = 3'b100;
	13'd3707: q = 3'b100;
	13'd3708: q = 3'b100;
	13'd3709: q = 3'b100;
	13'd3710: q = 3'b000;
	13'd3711: q = 3'b000;
	13'd3712: q = 3'b111;
	13'd3713: q = 3'b111;
	13'd3714: q = 3'b100;
	13'd3715: q = 3'b100;
	13'd3716: q = 3'b100;
	13'd3717: q = 3'b100;
	13'd3718: q = 3'b100;
	13'd3719: q = 3'b100;
	13'd3720: q = 3'b100;
	13'd3721: q = 3'b100;
	13'd3722: q = 3'b100;
	13'd3723: q = 3'b100;
	13'd3724: q = 3'b100;
	13'd3725: q = 3'b100;
	13'd3726: q = 3'b100;
	13'd3727: q = 3'b100;
	13'd3728: q = 3'b100;
	13'd3729: q = 3'b100;
	13'd3730: q = 3'b100;
	13'd3731: q = 3'b100;
	13'd3732: q = 3'b100;
	13'd3733: q = 3'b100;
	13'd3734: q = 3'b100;
	13'd3735: q = 3'b100;
	13'd3736: q = 3'b100;
	13'd3737: q = 3'b100;
	13'd3738: q = 3'b100;
	13'd3739: q = 3'b100;
	13'd3740: q = 3'b100;
	13'd3741: q = 3'b100;
	13'd3742: q = 3'b000;
	13'd3743: q = 3'b000;
	13'd3744: q = 3'b111;
	13'd3745: q = 3'b111;
	13'd3746: q = 3'b100;
	13'd3747: q = 3'b100;
	13'd3748: q = 3'b100;
	13'd3749: q = 3'b100;
	13'd3750: q = 3'b100;
	13'd3751: q = 3'b100;
	13'd3752: q = 3'b100;
	13'd3753: q = 3'b100;
	13'd3754: q = 3'b100;
	13'd3755: q = 3'b100;
	13'd3756: q = 3'b100;
	13'd3757: q = 3'b100;
	13'd3758: q = 3'b100;
	13'd3759: q = 3'b100;
	13'd3760: q = 3'b100;
	13'd3761: q = 3'b100;
	13'd3762: q = 3'b100;
	13'd3763: q = 3'b100;
	13'd3764: q = 3'b100;
	13'd3765: q = 3'b100;
	13'd3766: q = 3'b100;
	13'd3767: q = 3'b100;
	13'd3768: q = 3'b100;
	13'd3769: q = 3'b100;
	13'd3770: q = 3'b100;
	13'd3771: q = 3'b100;
	13'd3772: q = 3'b100;
	13'd3773: q = 3'b100;
	13'd3774: q = 3'b000;
	13'd3775: q = 3'b000;
	13'd3776: q = 3'b111;
	13'd3777: q = 3'b111;
	13'd3778: q = 3'b100;
	13'd3779: q = 3'b100;
	13'd3780: q = 3'b100;
	13'd3781: q = 3'b100;
	13'd3782: q = 3'b100;
	13'd3783: q = 3'b100;
	13'd3784: q = 3'b100;
	13'd3785: q = 3'b100;
	13'd3786: q = 3'b100;
	13'd3787: q = 3'b100;
	13'd3788: q = 3'b100;
	13'd3789: q = 3'b100;
	13'd3790: q = 3'b100;
	13'd3791: q = 3'b100;
	13'd3792: q = 3'b100;
	13'd3793: q = 3'b100;
	13'd3794: q = 3'b100;
	13'd3795: q = 3'b100;
	13'd3796: q = 3'b100;
	13'd3797: q = 3'b100;
	13'd3798: q = 3'b100;
	13'd3799: q = 3'b100;
	13'd3800: q = 3'b100;
	13'd3801: q = 3'b100;
	13'd3802: q = 3'b100;
	13'd3803: q = 3'b100;
	13'd3804: q = 3'b100;
	13'd3805: q = 3'b100;
	13'd3806: q = 3'b000;
	13'd3807: q = 3'b000;
	13'd3808: q = 3'b111;
	13'd3809: q = 3'b111;
	13'd3810: q = 3'b100;
	13'd3811: q = 3'b100;
	13'd3812: q = 3'b100;
	13'd3813: q = 3'b100;
	13'd3814: q = 3'b100;
	13'd3815: q = 3'b100;
	13'd3816: q = 3'b100;
	13'd3817: q = 3'b100;
	13'd3818: q = 3'b100;
	13'd3819: q = 3'b100;
	13'd3820: q = 3'b100;
	13'd3821: q = 3'b100;
	13'd3822: q = 3'b100;
	13'd3823: q = 3'b100;
	13'd3824: q = 3'b100;
	13'd3825: q = 3'b100;
	13'd3826: q = 3'b100;
	13'd3827: q = 3'b100;
	13'd3828: q = 3'b100;
	13'd3829: q = 3'b100;
	13'd3830: q = 3'b100;
	13'd3831: q = 3'b100;
	13'd3832: q = 3'b100;
	13'd3833: q = 3'b100;
	13'd3834: q = 3'b100;
	13'd3835: q = 3'b100;
	13'd3836: q = 3'b100;
	13'd3837: q = 3'b100;
	13'd3838: q = 3'b000;
	13'd3839: q = 3'b000;
	13'd3840: q = 3'b111;
	13'd3841: q = 3'b111;
	13'd3842: q = 3'b100;
	13'd3843: q = 3'b100;
	13'd3844: q = 3'b100;
	13'd3845: q = 3'b100;
	13'd3846: q = 3'b100;
	13'd3847: q = 3'b100;
	13'd3848: q = 3'b100;
	13'd3849: q = 3'b100;
	13'd3850: q = 3'b100;
	13'd3851: q = 3'b100;
	13'd3852: q = 3'b100;
	13'd3853: q = 3'b100;
	13'd3854: q = 3'b100;
	13'd3855: q = 3'b100;
	13'd3856: q = 3'b100;
	13'd3857: q = 3'b100;
	13'd3858: q = 3'b100;
	13'd3859: q = 3'b100;
	13'd3860: q = 3'b100;
	13'd3861: q = 3'b100;
	13'd3862: q = 3'b100;
	13'd3863: q = 3'b100;
	13'd3864: q = 3'b100;
	13'd3865: q = 3'b100;
	13'd3866: q = 3'b100;
	13'd3867: q = 3'b100;
	13'd3868: q = 3'b100;
	13'd3869: q = 3'b100;
	13'd3870: q = 3'b000;
	13'd3871: q = 3'b000;
	13'd3872: q = 3'b111;
	13'd3873: q = 3'b111;
	13'd3874: q = 3'b100;
	13'd3875: q = 3'b100;
	13'd3876: q = 3'b100;
	13'd3877: q = 3'b100;
	13'd3878: q = 3'b100;
	13'd3879: q = 3'b100;
	13'd3880: q = 3'b100;
	13'd3881: q = 3'b100;
	13'd3882: q = 3'b100;
	13'd3883: q = 3'b100;
	13'd3884: q = 3'b100;
	13'd3885: q = 3'b100;
	13'd3886: q = 3'b100;
	13'd3887: q = 3'b100;
	13'd3888: q = 3'b100;
	13'd3889: q = 3'b100;
	13'd3890: q = 3'b100;
	13'd3891: q = 3'b100;
	13'd3892: q = 3'b100;
	13'd3893: q = 3'b100;
	13'd3894: q = 3'b100;
	13'd3895: q = 3'b100;
	13'd3896: q = 3'b100;
	13'd3897: q = 3'b100;
	13'd3898: q = 3'b100;
	13'd3899: q = 3'b100;
	13'd3900: q = 3'b100;
	13'd3901: q = 3'b100;
	13'd3902: q = 3'b000;
	13'd3903: q = 3'b000;
	13'd3904: q = 3'b111;
	13'd3905: q = 3'b111;
	13'd3906: q = 3'b100;
	13'd3907: q = 3'b100;
	13'd3908: q = 3'b100;
	13'd3909: q = 3'b100;
	13'd3910: q = 3'b100;
	13'd3911: q = 3'b100;
	13'd3912: q = 3'b100;
	13'd3913: q = 3'b100;
	13'd3914: q = 3'b100;
	13'd3915: q = 3'b100;
	13'd3916: q = 3'b100;
	13'd3917: q = 3'b100;
	13'd3918: q = 3'b100;
	13'd3919: q = 3'b100;
	13'd3920: q = 3'b100;
	13'd3921: q = 3'b100;
	13'd3922: q = 3'b100;
	13'd3923: q = 3'b100;
	13'd3924: q = 3'b100;
	13'd3925: q = 3'b100;
	13'd3926: q = 3'b100;
	13'd3927: q = 3'b100;
	13'd3928: q = 3'b100;
	13'd3929: q = 3'b100;
	13'd3930: q = 3'b100;
	13'd3931: q = 3'b100;
	13'd3932: q = 3'b100;
	13'd3933: q = 3'b100;
	13'd3934: q = 3'b000;
	13'd3935: q = 3'b000;
	13'd3936: q = 3'b111;
	13'd3937: q = 3'b111;
	13'd3938: q = 3'b100;
	13'd3939: q = 3'b100;
	13'd3940: q = 3'b100;
	13'd3941: q = 3'b100;
	13'd3942: q = 3'b100;
	13'd3943: q = 3'b100;
	13'd3944: q = 3'b100;
	13'd3945: q = 3'b100;
	13'd3946: q = 3'b100;
	13'd3947: q = 3'b100;
	13'd3948: q = 3'b100;
	13'd3949: q = 3'b100;
	13'd3950: q = 3'b100;
	13'd3951: q = 3'b100;
	13'd3952: q = 3'b100;
	13'd3953: q = 3'b100;
	13'd3954: q = 3'b100;
	13'd3955: q = 3'b100;
	13'd3956: q = 3'b100;
	13'd3957: q = 3'b100;
	13'd3958: q = 3'b100;
	13'd3959: q = 3'b100;
	13'd3960: q = 3'b100;
	13'd3961: q = 3'b100;
	13'd3962: q = 3'b100;
	13'd3963: q = 3'b100;
	13'd3964: q = 3'b100;
	13'd3965: q = 3'b100;
	13'd3966: q = 3'b000;
	13'd3967: q = 3'b000;
	13'd3968: q = 3'b111;
	13'd3969: q = 3'b111;
	13'd3970: q = 3'b000;
	13'd3971: q = 3'b000;
	13'd3972: q = 3'b000;
	13'd3973: q = 3'b000;
	13'd3974: q = 3'b000;
	13'd3975: q = 3'b000;
	13'd3976: q = 3'b000;
	13'd3977: q = 3'b000;
	13'd3978: q = 3'b000;
	13'd3979: q = 3'b000;
	13'd3980: q = 3'b000;
	13'd3981: q = 3'b000;
	13'd3982: q = 3'b000;
	13'd3983: q = 3'b000;
	13'd3984: q = 3'b000;
	13'd3985: q = 3'b000;
	13'd3986: q = 3'b000;
	13'd3987: q = 3'b000;
	13'd3988: q = 3'b000;
	13'd3989: q = 3'b000;
	13'd3990: q = 3'b000;
	13'd3991: q = 3'b000;
	13'd3992: q = 3'b000;
	13'd3993: q = 3'b000;
	13'd3994: q = 3'b000;
	13'd3995: q = 3'b000;
	13'd3996: q = 3'b100;
	13'd3997: q = 3'b100;
	13'd3998: q = 3'b000;
	13'd3999: q = 3'b000;
	13'd4000: q = 3'b111;
	13'd4001: q = 3'b111;
	13'd4002: q = 3'b000;
	13'd4003: q = 3'b000;
	13'd4004: q = 3'b000;
	13'd4005: q = 3'b000;
	13'd4006: q = 3'b000;
	13'd4007: q = 3'b000;
	13'd4008: q = 3'b000;
	13'd4009: q = 3'b000;
	13'd4010: q = 3'b000;
	13'd4011: q = 3'b000;
	13'd4012: q = 3'b000;
	13'd4013: q = 3'b000;
	13'd4014: q = 3'b000;
	13'd4015: q = 3'b000;
	13'd4016: q = 3'b000;
	13'd4017: q = 3'b000;
	13'd4018: q = 3'b000;
	13'd4019: q = 3'b000;
	13'd4020: q = 3'b000;
	13'd4021: q = 3'b000;
	13'd4022: q = 3'b000;
	13'd4023: q = 3'b000;
	13'd4024: q = 3'b000;
	13'd4025: q = 3'b000;
	13'd4026: q = 3'b000;
	13'd4027: q = 3'b000;
	13'd4028: q = 3'b100;
	13'd4029: q = 3'b100;
	13'd4030: q = 3'b000;
	13'd4031: q = 3'b000;
	13'd4032: q = 3'b000;
	13'd4033: q = 3'b000;
	13'd4034: q = 3'b000;
	13'd4035: q = 3'b000;
	13'd4036: q = 3'b000;
	13'd4037: q = 3'b000;
	13'd4038: q = 3'b000;
	13'd4039: q = 3'b000;
	13'd4040: q = 3'b000;
	13'd4041: q = 3'b000;
	13'd4042: q = 3'b000;
	13'd4043: q = 3'b000;
	13'd4044: q = 3'b000;
	13'd4045: q = 3'b000;
	13'd4046: q = 3'b000;
	13'd4047: q = 3'b000;
	13'd4048: q = 3'b000;
	13'd4049: q = 3'b000;
	13'd4050: q = 3'b000;
	13'd4051: q = 3'b000;
	13'd4052: q = 3'b000;
	13'd4053: q = 3'b000;
	13'd4054: q = 3'b000;
	13'd4055: q = 3'b000;
	13'd4056: q = 3'b000;
	13'd4057: q = 3'b000;
	13'd4058: q = 3'b000;
	13'd4059: q = 3'b000;
	13'd4060: q = 3'b000;
	13'd4061: q = 3'b000;
	13'd4062: q = 3'b000;
	13'd4063: q = 3'b000;
	13'd4064: q = 3'b000;
	13'd4065: q = 3'b000;
	13'd4066: q = 3'b000;
	13'd4067: q = 3'b000;
	13'd4068: q = 3'b000;
	13'd4069: q = 3'b000;
	13'd4070: q = 3'b000;
	13'd4071: q = 3'b000;
	13'd4072: q = 3'b000;
	13'd4073: q = 3'b000;
	13'd4074: q = 3'b000;
	13'd4075: q = 3'b000;
	13'd4076: q = 3'b000;
	13'd4077: q = 3'b000;
	13'd4078: q = 3'b000;
	13'd4079: q = 3'b000;
	13'd4080: q = 3'b000;
	13'd4081: q = 3'b000;
	13'd4082: q = 3'b000;
	13'd4083: q = 3'b000;
	13'd4084: q = 3'b000;
	13'd4085: q = 3'b000;
	13'd4086: q = 3'b000;
	13'd4087: q = 3'b000;
	13'd4088: q = 3'b000;
	13'd4089: q = 3'b000;
	13'd4090: q = 3'b000;
	13'd4091: q = 3'b000;
	13'd4092: q = 3'b000;
	13'd4093: q = 3'b000;
	13'd4094: q = 3'b000;
	13'd4095: q = 3'b000;
	13'd4096: q = 3'b000;
	13'd4097: q = 3'b000;
	13'd4098: q = 3'b000;
	13'd4099: q = 3'b000;
	13'd4100: q = 3'b000;
	13'd4101: q = 3'b000;
	13'd4102: q = 3'b000;
	13'd4103: q = 3'b000;
	13'd4104: q = 3'b000;
	13'd4105: q = 3'b000;
	13'd4106: q = 3'b000;
	13'd4107: q = 3'b000;
	13'd4108: q = 3'b000;
	13'd4109: q = 3'b000;
	13'd4110: q = 3'b000;
	13'd4111: q = 3'b000;
	13'd4112: q = 3'b000;
	13'd4113: q = 3'b000;
	13'd4114: q = 3'b000;
	13'd4115: q = 3'b000;
	13'd4116: q = 3'b000;
	13'd4117: q = 3'b000;
	13'd4118: q = 3'b000;
	13'd4119: q = 3'b000;
	13'd4120: q = 3'b000;
	13'd4121: q = 3'b000;
	13'd4122: q = 3'b000;
	13'd4123: q = 3'b000;
	13'd4124: q = 3'b000;
	13'd4125: q = 3'b000;
	13'd4126: q = 3'b000;
	13'd4127: q = 3'b000;
	13'd4128: q = 3'b000;
	13'd4129: q = 3'b000;
	13'd4130: q = 3'b000;
	13'd4131: q = 3'b000;
	13'd4132: q = 3'b000;
	13'd4133: q = 3'b000;
	13'd4134: q = 3'b000;
	13'd4135: q = 3'b000;
	13'd4136: q = 3'b000;
	13'd4137: q = 3'b000;
	13'd4138: q = 3'b000;
	13'd4139: q = 3'b000;
	13'd4140: q = 3'b000;
	13'd4141: q = 3'b000;
	13'd4142: q = 3'b000;
	13'd4143: q = 3'b000;
	13'd4144: q = 3'b000;
	13'd4145: q = 3'b000;
	13'd4146: q = 3'b000;
	13'd4147: q = 3'b000;
	13'd4148: q = 3'b000;
	13'd4149: q = 3'b000;
	13'd4150: q = 3'b000;
	13'd4151: q = 3'b000;
	13'd4152: q = 3'b000;
	13'd4153: q = 3'b000;
	13'd4154: q = 3'b000;
	13'd4155: q = 3'b000;
	13'd4156: q = 3'b000;
	13'd4157: q = 3'b000;
	13'd4158: q = 3'b000;
	13'd4159: q = 3'b000;
	13'd4160: q = 3'b000;
	13'd4161: q = 3'b000;
	13'd4162: q = 3'b111;
	13'd4163: q = 3'b111;
	13'd4164: q = 3'b111;
	13'd4165: q = 3'b111;
	13'd4166: q = 3'b111;
	13'd4167: q = 3'b111;
	13'd4168: q = 3'b111;
	13'd4169: q = 3'b111;
	13'd4170: q = 3'b111;
	13'd4171: q = 3'b111;
	13'd4172: q = 3'b111;
	13'd4173: q = 3'b111;
	13'd4174: q = 3'b111;
	13'd4175: q = 3'b111;
	13'd4176: q = 3'b111;
	13'd4177: q = 3'b111;
	13'd4178: q = 3'b111;
	13'd4179: q = 3'b111;
	13'd4180: q = 3'b111;
	13'd4181: q = 3'b111;
	13'd4182: q = 3'b111;
	13'd4183: q = 3'b111;
	13'd4184: q = 3'b111;
	13'd4185: q = 3'b111;
	13'd4186: q = 3'b111;
	13'd4187: q = 3'b111;
	13'd4188: q = 3'b111;
	13'd4189: q = 3'b111;
	13'd4190: q = 3'b000;
	13'd4191: q = 3'b000;
	13'd4192: q = 3'b000;
	13'd4193: q = 3'b000;
	13'd4194: q = 3'b111;
	13'd4195: q = 3'b111;
	13'd4196: q = 3'b111;
	13'd4197: q = 3'b111;
	13'd4198: q = 3'b111;
	13'd4199: q = 3'b111;
	13'd4200: q = 3'b111;
	13'd4201: q = 3'b111;
	13'd4202: q = 3'b111;
	13'd4203: q = 3'b111;
	13'd4204: q = 3'b111;
	13'd4205: q = 3'b111;
	13'd4206: q = 3'b111;
	13'd4207: q = 3'b111;
	13'd4208: q = 3'b111;
	13'd4209: q = 3'b111;
	13'd4210: q = 3'b111;
	13'd4211: q = 3'b111;
	13'd4212: q = 3'b111;
	13'd4213: q = 3'b111;
	13'd4214: q = 3'b111;
	13'd4215: q = 3'b111;
	13'd4216: q = 3'b111;
	13'd4217: q = 3'b111;
	13'd4218: q = 3'b111;
	13'd4219: q = 3'b111;
	13'd4220: q = 3'b111;
	13'd4221: q = 3'b111;
	13'd4222: q = 3'b000;
	13'd4223: q = 3'b000;
	13'd4224: q = 3'b111;
	13'd4225: q = 3'b111;
	13'd4226: q = 3'b100;
	13'd4227: q = 3'b100;
	13'd4228: q = 3'b100;
	13'd4229: q = 3'b100;
	13'd4230: q = 3'b100;
	13'd4231: q = 3'b100;
	13'd4232: q = 3'b100;
	13'd4233: q = 3'b100;
	13'd4234: q = 3'b100;
	13'd4235: q = 3'b100;
	13'd4236: q = 3'b100;
	13'd4237: q = 3'b100;
	13'd4238: q = 3'b100;
	13'd4239: q = 3'b100;
	13'd4240: q = 3'b100;
	13'd4241: q = 3'b100;
	13'd4242: q = 3'b100;
	13'd4243: q = 3'b100;
	13'd4244: q = 3'b100;
	13'd4245: q = 3'b100;
	13'd4246: q = 3'b100;
	13'd4247: q = 3'b100;
	13'd4248: q = 3'b100;
	13'd4249: q = 3'b100;
	13'd4250: q = 3'b100;
	13'd4251: q = 3'b100;
	13'd4252: q = 3'b100;
	13'd4253: q = 3'b100;
	13'd4254: q = 3'b000;
	13'd4255: q = 3'b000;
	13'd4256: q = 3'b111;
	13'd4257: q = 3'b111;
	13'd4258: q = 3'b100;
	13'd4259: q = 3'b100;
	13'd4260: q = 3'b100;
	13'd4261: q = 3'b100;
	13'd4262: q = 3'b100;
	13'd4263: q = 3'b100;
	13'd4264: q = 3'b100;
	13'd4265: q = 3'b100;
	13'd4266: q = 3'b100;
	13'd4267: q = 3'b100;
	13'd4268: q = 3'b100;
	13'd4269: q = 3'b100;
	13'd4270: q = 3'b100;
	13'd4271: q = 3'b100;
	13'd4272: q = 3'b100;
	13'd4273: q = 3'b100;
	13'd4274: q = 3'b100;
	13'd4275: q = 3'b100;
	13'd4276: q = 3'b100;
	13'd4277: q = 3'b100;
	13'd4278: q = 3'b100;
	13'd4279: q = 3'b100;
	13'd4280: q = 3'b100;
	13'd4281: q = 3'b100;
	13'd4282: q = 3'b100;
	13'd4283: q = 3'b100;
	13'd4284: q = 3'b100;
	13'd4285: q = 3'b100;
	13'd4286: q = 3'b000;
	13'd4287: q = 3'b000;
	13'd4288: q = 3'b111;
	13'd4289: q = 3'b111;
	13'd4290: q = 3'b100;
	13'd4291: q = 3'b100;
	13'd4292: q = 3'b100;
	13'd4293: q = 3'b100;
	13'd4294: q = 3'b100;
	13'd4295: q = 3'b100;
	13'd4296: q = 3'b100;
	13'd4297: q = 3'b100;
	13'd4298: q = 3'b100;
	13'd4299: q = 3'b100;
	13'd4300: q = 3'b100;
	13'd4301: q = 3'b100;
	13'd4302: q = 3'b100;
	13'd4303: q = 3'b100;
	13'd4304: q = 3'b100;
	13'd4305: q = 3'b100;
	13'd4306: q = 3'b100;
	13'd4307: q = 3'b100;
	13'd4308: q = 3'b100;
	13'd4309: q = 3'b100;
	13'd4310: q = 3'b100;
	13'd4311: q = 3'b100;
	13'd4312: q = 3'b100;
	13'd4313: q = 3'b100;
	13'd4314: q = 3'b100;
	13'd4315: q = 3'b100;
	13'd4316: q = 3'b100;
	13'd4317: q = 3'b100;
	13'd4318: q = 3'b000;
	13'd4319: q = 3'b000;
	13'd4320: q = 3'b111;
	13'd4321: q = 3'b111;
	13'd4322: q = 3'b100;
	13'd4323: q = 3'b100;
	13'd4324: q = 3'b100;
	13'd4325: q = 3'b100;
	13'd4326: q = 3'b100;
	13'd4327: q = 3'b100;
	13'd4328: q = 3'b100;
	13'd4329: q = 3'b100;
	13'd4330: q = 3'b100;
	13'd4331: q = 3'b100;
	13'd4332: q = 3'b100;
	13'd4333: q = 3'b100;
	13'd4334: q = 3'b100;
	13'd4335: q = 3'b100;
	13'd4336: q = 3'b100;
	13'd4337: q = 3'b100;
	13'd4338: q = 3'b100;
	13'd4339: q = 3'b100;
	13'd4340: q = 3'b100;
	13'd4341: q = 3'b100;
	13'd4342: q = 3'b100;
	13'd4343: q = 3'b100;
	13'd4344: q = 3'b100;
	13'd4345: q = 3'b100;
	13'd4346: q = 3'b100;
	13'd4347: q = 3'b100;
	13'd4348: q = 3'b100;
	13'd4349: q = 3'b100;
	13'd4350: q = 3'b000;
	13'd4351: q = 3'b000;
	13'd4352: q = 3'b111;
	13'd4353: q = 3'b111;
	13'd4354: q = 3'b100;
	13'd4355: q = 3'b100;
	13'd4356: q = 3'b100;
	13'd4357: q = 3'b100;
	13'd4358: q = 3'b100;
	13'd4359: q = 3'b100;
	13'd4360: q = 3'b100;
	13'd4361: q = 3'b100;
	13'd4362: q = 3'b100;
	13'd4363: q = 3'b100;
	13'd4364: q = 3'b100;
	13'd4365: q = 3'b100;
	13'd4366: q = 3'b100;
	13'd4367: q = 3'b100;
	13'd4368: q = 3'b100;
	13'd4369: q = 3'b100;
	13'd4370: q = 3'b100;
	13'd4371: q = 3'b100;
	13'd4372: q = 3'b100;
	13'd4373: q = 3'b100;
	13'd4374: q = 3'b100;
	13'd4375: q = 3'b100;
	13'd4376: q = 3'b100;
	13'd4377: q = 3'b100;
	13'd4378: q = 3'b100;
	13'd4379: q = 3'b100;
	13'd4380: q = 3'b100;
	13'd4381: q = 3'b100;
	13'd4382: q = 3'b000;
	13'd4383: q = 3'b000;
	13'd4384: q = 3'b111;
	13'd4385: q = 3'b111;
	13'd4386: q = 3'b100;
	13'd4387: q = 3'b100;
	13'd4388: q = 3'b100;
	13'd4389: q = 3'b100;
	13'd4390: q = 3'b100;
	13'd4391: q = 3'b100;
	13'd4392: q = 3'b100;
	13'd4393: q = 3'b100;
	13'd4394: q = 3'b100;
	13'd4395: q = 3'b100;
	13'd4396: q = 3'b100;
	13'd4397: q = 3'b100;
	13'd4398: q = 3'b100;
	13'd4399: q = 3'b100;
	13'd4400: q = 3'b100;
	13'd4401: q = 3'b100;
	13'd4402: q = 3'b100;
	13'd4403: q = 3'b100;
	13'd4404: q = 3'b100;
	13'd4405: q = 3'b100;
	13'd4406: q = 3'b100;
	13'd4407: q = 3'b100;
	13'd4408: q = 3'b100;
	13'd4409: q = 3'b100;
	13'd4410: q = 3'b100;
	13'd4411: q = 3'b100;
	13'd4412: q = 3'b100;
	13'd4413: q = 3'b100;
	13'd4414: q = 3'b000;
	13'd4415: q = 3'b000;
	13'd4416: q = 3'b000;
	13'd4417: q = 3'b000;
	13'd4418: q = 3'b000;
	13'd4419: q = 3'b000;
	13'd4420: q = 3'b000;
	13'd4421: q = 3'b000;
	13'd4422: q = 3'b000;
	13'd4423: q = 3'b000;
	13'd4424: q = 3'b000;
	13'd4425: q = 3'b000;
	13'd4426: q = 3'b000;
	13'd4427: q = 3'b000;
	13'd4428: q = 3'b000;
	13'd4429: q = 3'b000;
	13'd4430: q = 3'b000;
	13'd4431: q = 3'b000;
	13'd4432: q = 3'b000;
	13'd4433: q = 3'b000;
	13'd4434: q = 3'b000;
	13'd4435: q = 3'b000;
	13'd4436: q = 3'b000;
	13'd4437: q = 3'b000;
	13'd4438: q = 3'b000;
	13'd4439: q = 3'b000;
	13'd4440: q = 3'b000;
	13'd4441: q = 3'b000;
	13'd4442: q = 3'b000;
	13'd4443: q = 3'b000;
	13'd4444: q = 3'b000;
	13'd4445: q = 3'b000;
	13'd4446: q = 3'b000;
	13'd4447: q = 3'b000;
	13'd4448: q = 3'b000;
	13'd4449: q = 3'b000;
	13'd4450: q = 3'b000;
	13'd4451: q = 3'b000;
	13'd4452: q = 3'b000;
	13'd4453: q = 3'b000;
	13'd4454: q = 3'b000;
	13'd4455: q = 3'b000;
	13'd4456: q = 3'b000;
	13'd4457: q = 3'b000;
	13'd4458: q = 3'b000;
	13'd4459: q = 3'b000;
	13'd4460: q = 3'b000;
	13'd4461: q = 3'b000;
	13'd4462: q = 3'b000;
	13'd4463: q = 3'b000;
	13'd4464: q = 3'b000;
	13'd4465: q = 3'b000;
	13'd4466: q = 3'b000;
	13'd4467: q = 3'b000;
	13'd4468: q = 3'b000;
	13'd4469: q = 3'b000;
	13'd4470: q = 3'b000;
	13'd4471: q = 3'b000;
	13'd4472: q = 3'b000;
	13'd4473: q = 3'b000;
	13'd4474: q = 3'b000;
	13'd4475: q = 3'b000;
	13'd4476: q = 3'b000;
	13'd4477: q = 3'b000;
	13'd4478: q = 3'b000;
	13'd4479: q = 3'b000;
	13'd4480: q = 3'b111;
	13'd4481: q = 3'b111;
	13'd4482: q = 3'b111;
	13'd4483: q = 3'b111;
	13'd4484: q = 3'b111;
	13'd4485: q = 3'b111;
	13'd4486: q = 3'b111;
	13'd4487: q = 3'b111;
	13'd4488: q = 3'b111;
	13'd4489: q = 3'b111;
	13'd4490: q = 3'b000;
	13'd4491: q = 3'b000;
	13'd4492: q = 3'b000;
	13'd4493: q = 3'b000;
	13'd4494: q = 3'b111;
	13'd4495: q = 3'b111;
	13'd4496: q = 3'b111;
	13'd4497: q = 3'b111;
	13'd4498: q = 3'b111;
	13'd4499: q = 3'b111;
	13'd4500: q = 3'b111;
	13'd4501: q = 3'b111;
	13'd4502: q = 3'b111;
	13'd4503: q = 3'b111;
	13'd4504: q = 3'b111;
	13'd4505: q = 3'b111;
	13'd4506: q = 3'b111;
	13'd4507: q = 3'b111;
	13'd4508: q = 3'b111;
	13'd4509: q = 3'b111;
	13'd4510: q = 3'b111;
	13'd4511: q = 3'b111;
	13'd4512: q = 3'b111;
	13'd4513: q = 3'b111;
	13'd4514: q = 3'b111;
	13'd4515: q = 3'b111;
	13'd4516: q = 3'b111;
	13'd4517: q = 3'b111;
	13'd4518: q = 3'b111;
	13'd4519: q = 3'b111;
	13'd4520: q = 3'b111;
	13'd4521: q = 3'b111;
	13'd4522: q = 3'b000;
	13'd4523: q = 3'b000;
	13'd4524: q = 3'b000;
	13'd4525: q = 3'b000;
	13'd4526: q = 3'b111;
	13'd4527: q = 3'b111;
	13'd4528: q = 3'b111;
	13'd4529: q = 3'b111;
	13'd4530: q = 3'b111;
	13'd4531: q = 3'b111;
	13'd4532: q = 3'b111;
	13'd4533: q = 3'b111;
	13'd4534: q = 3'b111;
	13'd4535: q = 3'b111;
	13'd4536: q = 3'b111;
	13'd4537: q = 3'b111;
	13'd4538: q = 3'b111;
	13'd4539: q = 3'b111;
	13'd4540: q = 3'b111;
	13'd4541: q = 3'b111;
	13'd4542: q = 3'b111;
	13'd4543: q = 3'b111;
	13'd4544: q = 3'b100;
	13'd4545: q = 3'b100;
	13'd4546: q = 3'b100;
	13'd4547: q = 3'b100;
	13'd4548: q = 3'b100;
	13'd4549: q = 3'b100;
	13'd4550: q = 3'b100;
	13'd4551: q = 3'b100;
	13'd4552: q = 3'b100;
	13'd4553: q = 3'b100;
	13'd4554: q = 3'b000;
	13'd4555: q = 3'b000;
	13'd4556: q = 3'b111;
	13'd4557: q = 3'b111;
	13'd4558: q = 3'b100;
	13'd4559: q = 3'b100;
	13'd4560: q = 3'b100;
	13'd4561: q = 3'b100;
	13'd4562: q = 3'b100;
	13'd4563: q = 3'b100;
	13'd4564: q = 3'b100;
	13'd4565: q = 3'b100;
	13'd4566: q = 3'b100;
	13'd4567: q = 3'b100;
	13'd4568: q = 3'b100;
	13'd4569: q = 3'b100;
	13'd4570: q = 3'b100;
	13'd4571: q = 3'b100;
	13'd4572: q = 3'b100;
	13'd4573: q = 3'b100;
	13'd4574: q = 3'b100;
	13'd4575: q = 3'b100;
	13'd4576: q = 3'b100;
	13'd4577: q = 3'b100;
	13'd4578: q = 3'b100;
	13'd4579: q = 3'b100;
	13'd4580: q = 3'b100;
	13'd4581: q = 3'b100;
	13'd4582: q = 3'b100;
	13'd4583: q = 3'b100;
	13'd4584: q = 3'b100;
	13'd4585: q = 3'b100;
	13'd4586: q = 3'b000;
	13'd4587: q = 3'b000;
	13'd4588: q = 3'b111;
	13'd4589: q = 3'b111;
	13'd4590: q = 3'b100;
	13'd4591: q = 3'b100;
	13'd4592: q = 3'b100;
	13'd4593: q = 3'b100;
	13'd4594: q = 3'b100;
	13'd4595: q = 3'b100;
	13'd4596: q = 3'b100;
	13'd4597: q = 3'b100;
	13'd4598: q = 3'b100;
	13'd4599: q = 3'b100;
	13'd4600: q = 3'b100;
	13'd4601: q = 3'b100;
	13'd4602: q = 3'b100;
	13'd4603: q = 3'b100;
	13'd4604: q = 3'b100;
	13'd4605: q = 3'b100;
	13'd4606: q = 3'b100;
	13'd4607: q = 3'b100;
	13'd4608: q = 3'b100;
	13'd4609: q = 3'b100;
	13'd4610: q = 3'b100;
	13'd4611: q = 3'b100;
	13'd4612: q = 3'b100;
	13'd4613: q = 3'b100;
	13'd4614: q = 3'b100;
	13'd4615: q = 3'b100;
	13'd4616: q = 3'b100;
	13'd4617: q = 3'b100;
	13'd4618: q = 3'b000;
	13'd4619: q = 3'b000;
	13'd4620: q = 3'b111;
	13'd4621: q = 3'b111;
	13'd4622: q = 3'b100;
	13'd4623: q = 3'b100;
	13'd4624: q = 3'b100;
	13'd4625: q = 3'b100;
	13'd4626: q = 3'b100;
	13'd4627: q = 3'b100;
	13'd4628: q = 3'b100;
	13'd4629: q = 3'b100;
	13'd4630: q = 3'b100;
	13'd4631: q = 3'b100;
	13'd4632: q = 3'b100;
	13'd4633: q = 3'b100;
	13'd4634: q = 3'b100;
	13'd4635: q = 3'b100;
	13'd4636: q = 3'b100;
	13'd4637: q = 3'b100;
	13'd4638: q = 3'b100;
	13'd4639: q = 3'b100;
	13'd4640: q = 3'b100;
	13'd4641: q = 3'b100;
	13'd4642: q = 3'b100;
	13'd4643: q = 3'b100;
	13'd4644: q = 3'b100;
	13'd4645: q = 3'b100;
	13'd4646: q = 3'b100;
	13'd4647: q = 3'b100;
	13'd4648: q = 3'b100;
	13'd4649: q = 3'b100;
	13'd4650: q = 3'b000;
	13'd4651: q = 3'b000;
	13'd4652: q = 3'b111;
	13'd4653: q = 3'b111;
	13'd4654: q = 3'b100;
	13'd4655: q = 3'b100;
	13'd4656: q = 3'b100;
	13'd4657: q = 3'b100;
	13'd4658: q = 3'b100;
	13'd4659: q = 3'b100;
	13'd4660: q = 3'b100;
	13'd4661: q = 3'b100;
	13'd4662: q = 3'b100;
	13'd4663: q = 3'b100;
	13'd4664: q = 3'b100;
	13'd4665: q = 3'b100;
	13'd4666: q = 3'b100;
	13'd4667: q = 3'b100;
	13'd4668: q = 3'b100;
	13'd4669: q = 3'b100;
	13'd4670: q = 3'b100;
	13'd4671: q = 3'b100;
	13'd4672: q = 3'b100;
	13'd4673: q = 3'b100;
	13'd4674: q = 3'b100;
	13'd4675: q = 3'b100;
	13'd4676: q = 3'b100;
	13'd4677: q = 3'b100;
	13'd4678: q = 3'b100;
	13'd4679: q = 3'b100;
	13'd4680: q = 3'b100;
	13'd4681: q = 3'b100;
	13'd4682: q = 3'b000;
	13'd4683: q = 3'b000;
	13'd4684: q = 3'b111;
	13'd4685: q = 3'b111;
	13'd4686: q = 3'b100;
	13'd4687: q = 3'b100;
	13'd4688: q = 3'b100;
	13'd4689: q = 3'b100;
	13'd4690: q = 3'b100;
	13'd4691: q = 3'b100;
	13'd4692: q = 3'b100;
	13'd4693: q = 3'b100;
	13'd4694: q = 3'b100;
	13'd4695: q = 3'b100;
	13'd4696: q = 3'b100;
	13'd4697: q = 3'b100;
	13'd4698: q = 3'b100;
	13'd4699: q = 3'b100;
	13'd4700: q = 3'b100;
	13'd4701: q = 3'b100;
	13'd4702: q = 3'b100;
	13'd4703: q = 3'b100;
	13'd4704: q = 3'b100;
	13'd4705: q = 3'b100;
	13'd4706: q = 3'b100;
	13'd4707: q = 3'b100;
	13'd4708: q = 3'b100;
	13'd4709: q = 3'b100;
	13'd4710: q = 3'b100;
	13'd4711: q = 3'b100;
	13'd4712: q = 3'b100;
	13'd4713: q = 3'b100;
	13'd4714: q = 3'b000;
	13'd4715: q = 3'b000;
	13'd4716: q = 3'b111;
	13'd4717: q = 3'b111;
	13'd4718: q = 3'b100;
	13'd4719: q = 3'b100;
	13'd4720: q = 3'b100;
	13'd4721: q = 3'b100;
	13'd4722: q = 3'b100;
	13'd4723: q = 3'b100;
	13'd4724: q = 3'b100;
	13'd4725: q = 3'b100;
	13'd4726: q = 3'b100;
	13'd4727: q = 3'b100;
	13'd4728: q = 3'b100;
	13'd4729: q = 3'b100;
	13'd4730: q = 3'b100;
	13'd4731: q = 3'b100;
	13'd4732: q = 3'b100;
	13'd4733: q = 3'b100;
	13'd4734: q = 3'b100;
	13'd4735: q = 3'b100;
	13'd4736: q = 3'b000;
	13'd4737: q = 3'b000;
	13'd4738: q = 3'b000;
	13'd4739: q = 3'b000;
	13'd4740: q = 3'b000;
	13'd4741: q = 3'b000;
	13'd4742: q = 3'b000;
	13'd4743: q = 3'b000;
	13'd4744: q = 3'b000;
	13'd4745: q = 3'b000;
	13'd4746: q = 3'b000;
	13'd4747: q = 3'b000;
	13'd4748: q = 3'b000;
	13'd4749: q = 3'b000;
	13'd4750: q = 3'b000;
	13'd4751: q = 3'b000;
	13'd4752: q = 3'b000;
	13'd4753: q = 3'b000;
	13'd4754: q = 3'b000;
	13'd4755: q = 3'b000;
	13'd4756: q = 3'b000;
	13'd4757: q = 3'b000;
	13'd4758: q = 3'b000;
	13'd4759: q = 3'b000;
	13'd4760: q = 3'b000;
	13'd4761: q = 3'b000;
	13'd4762: q = 3'b000;
	13'd4763: q = 3'b000;
	13'd4764: q = 3'b000;
	13'd4765: q = 3'b000;
	13'd4766: q = 3'b000;
	13'd4767: q = 3'b000;
	13'd4768: q = 3'b000;
	13'd4769: q = 3'b000;
	13'd4770: q = 3'b000;
	13'd4771: q = 3'b000;
	13'd4772: q = 3'b000;
	13'd4773: q = 3'b000;
	13'd4774: q = 3'b000;
	13'd4775: q = 3'b000;
	13'd4776: q = 3'b000;
	13'd4777: q = 3'b000;
	13'd4778: q = 3'b000;
	13'd4779: q = 3'b000;
	13'd4780: q = 3'b000;
	13'd4781: q = 3'b000;
	13'd4782: q = 3'b000;
	13'd4783: q = 3'b000;
	13'd4784: q = 3'b000;
	13'd4785: q = 3'b000;
	13'd4786: q = 3'b000;
	13'd4787: q = 3'b000;
	13'd4788: q = 3'b000;
	13'd4789: q = 3'b000;
	13'd4790: q = 3'b000;
	13'd4791: q = 3'b000;
	13'd4792: q = 3'b000;
	13'd4793: q = 3'b000;
	13'd4794: q = 3'b000;
	13'd4795: q = 3'b000;
	13'd4796: q = 3'b000;
	13'd4797: q = 3'b000;
	13'd4798: q = 3'b000;
	13'd4799: q = 3'b000;
	13'd4800: q = 3'b111;
	13'd4801: q = 3'b111;
	13'd4802: q = 3'b111;
	13'd4803: q = 3'b111;
	13'd4804: q = 3'b111;
	13'd4805: q = 3'b111;
	13'd4806: q = 3'b111;
	13'd4807: q = 3'b111;
	13'd4808: q = 3'b111;
	13'd4809: q = 3'b111;
	13'd4810: q = 3'b111;
	13'd4811: q = 3'b111;
	13'd4812: q = 3'b111;
	13'd4813: q = 3'b111;
	13'd4814: q = 3'b111;
	13'd4815: q = 3'b111;
	13'd4816: q = 3'b111;
	13'd4817: q = 3'b111;
	13'd4818: q = 3'b000;
	13'd4819: q = 3'b000;
	13'd4820: q = 3'b000;
	13'd4821: q = 3'b000;
	13'd4822: q = 3'b111;
	13'd4823: q = 3'b111;
	13'd4824: q = 3'b111;
	13'd4825: q = 3'b111;
	13'd4826: q = 3'b111;
	13'd4827: q = 3'b111;
	13'd4828: q = 3'b111;
	13'd4829: q = 3'b111;
	13'd4830: q = 3'b111;
	13'd4831: q = 3'b111;
	13'd4832: q = 3'b111;
	13'd4833: q = 3'b111;
	13'd4834: q = 3'b111;
	13'd4835: q = 3'b111;
	13'd4836: q = 3'b111;
	13'd4837: q = 3'b111;
	13'd4838: q = 3'b111;
	13'd4839: q = 3'b111;
	13'd4840: q = 3'b111;
	13'd4841: q = 3'b111;
	13'd4842: q = 3'b111;
	13'd4843: q = 3'b111;
	13'd4844: q = 3'b111;
	13'd4845: q = 3'b111;
	13'd4846: q = 3'b111;
	13'd4847: q = 3'b111;
	13'd4848: q = 3'b111;
	13'd4849: q = 3'b111;
	13'd4850: q = 3'b000;
	13'd4851: q = 3'b000;
	13'd4852: q = 3'b000;
	13'd4853: q = 3'b000;
	13'd4854: q = 3'b111;
	13'd4855: q = 3'b111;
	13'd4856: q = 3'b111;
	13'd4857: q = 3'b111;
	13'd4858: q = 3'b111;
	13'd4859: q = 3'b111;
	13'd4860: q = 3'b111;
	13'd4861: q = 3'b111;
	13'd4862: q = 3'b111;
	13'd4863: q = 3'b111;
	13'd4864: q = 3'b100;
	13'd4865: q = 3'b100;
	13'd4866: q = 3'b100;
	13'd4867: q = 3'b100;
	13'd4868: q = 3'b100;
	13'd4869: q = 3'b100;
	13'd4870: q = 3'b100;
	13'd4871: q = 3'b100;
	13'd4872: q = 3'b100;
	13'd4873: q = 3'b100;
	13'd4874: q = 3'b100;
	13'd4875: q = 3'b100;
	13'd4876: q = 3'b100;
	13'd4877: q = 3'b100;
	13'd4878: q = 3'b100;
	13'd4879: q = 3'b100;
	13'd4880: q = 3'b100;
	13'd4881: q = 3'b100;
	13'd4882: q = 3'b000;
	13'd4883: q = 3'b000;
	13'd4884: q = 3'b111;
	13'd4885: q = 3'b111;
	13'd4886: q = 3'b100;
	13'd4887: q = 3'b100;
	13'd4888: q = 3'b100;
	13'd4889: q = 3'b100;
	13'd4890: q = 3'b100;
	13'd4891: q = 3'b100;
	13'd4892: q = 3'b100;
	13'd4893: q = 3'b100;
	13'd4894: q = 3'b100;
	13'd4895: q = 3'b100;
	13'd4896: q = 3'b100;
	13'd4897: q = 3'b100;
	13'd4898: q = 3'b100;
	13'd4899: q = 3'b100;
	13'd4900: q = 3'b100;
	13'd4901: q = 3'b100;
	13'd4902: q = 3'b100;
	13'd4903: q = 3'b100;
	13'd4904: q = 3'b100;
	13'd4905: q = 3'b100;
	13'd4906: q = 3'b100;
	13'd4907: q = 3'b100;
	13'd4908: q = 3'b100;
	13'd4909: q = 3'b100;
	13'd4910: q = 3'b100;
	13'd4911: q = 3'b100;
	13'd4912: q = 3'b100;
	13'd4913: q = 3'b100;
	13'd4914: q = 3'b000;
	13'd4915: q = 3'b000;
	13'd4916: q = 3'b111;
	13'd4917: q = 3'b111;
	13'd4918: q = 3'b100;
	13'd4919: q = 3'b100;
	13'd4920: q = 3'b100;
	13'd4921: q = 3'b100;
	13'd4922: q = 3'b100;
	13'd4923: q = 3'b100;
	13'd4924: q = 3'b100;
	13'd4925: q = 3'b100;
	13'd4926: q = 3'b100;
	13'd4927: q = 3'b100;
	13'd4928: q = 3'b100;
	13'd4929: q = 3'b100;
	13'd4930: q = 3'b100;
	13'd4931: q = 3'b100;
	13'd4932: q = 3'b100;
	13'd4933: q = 3'b100;
	13'd4934: q = 3'b100;
	13'd4935: q = 3'b100;
	13'd4936: q = 3'b100;
	13'd4937: q = 3'b100;
	13'd4938: q = 3'b100;
	13'd4939: q = 3'b100;
	13'd4940: q = 3'b100;
	13'd4941: q = 3'b100;
	13'd4942: q = 3'b100;
	13'd4943: q = 3'b100;
	13'd4944: q = 3'b100;
	13'd4945: q = 3'b100;
	13'd4946: q = 3'b000;
	13'd4947: q = 3'b000;
	13'd4948: q = 3'b111;
	13'd4949: q = 3'b111;
	13'd4950: q = 3'b100;
	13'd4951: q = 3'b100;
	13'd4952: q = 3'b100;
	13'd4953: q = 3'b100;
	13'd4954: q = 3'b100;
	13'd4955: q = 3'b100;
	13'd4956: q = 3'b100;
	13'd4957: q = 3'b100;
	13'd4958: q = 3'b100;
	13'd4959: q = 3'b100;
	13'd4960: q = 3'b100;
	13'd4961: q = 3'b100;
	13'd4962: q = 3'b100;
	13'd4963: q = 3'b100;
	13'd4964: q = 3'b100;
	13'd4965: q = 3'b100;
	13'd4966: q = 3'b100;
	13'd4967: q = 3'b100;
	13'd4968: q = 3'b100;
	13'd4969: q = 3'b100;
	13'd4970: q = 3'b100;
	13'd4971: q = 3'b100;
	13'd4972: q = 3'b100;
	13'd4973: q = 3'b100;
	13'd4974: q = 3'b100;
	13'd4975: q = 3'b100;
	13'd4976: q = 3'b100;
	13'd4977: q = 3'b100;
	13'd4978: q = 3'b000;
	13'd4979: q = 3'b000;
	13'd4980: q = 3'b111;
	13'd4981: q = 3'b111;
	13'd4982: q = 3'b100;
	13'd4983: q = 3'b100;
	13'd4984: q = 3'b100;
	13'd4985: q = 3'b100;
	13'd4986: q = 3'b100;
	13'd4987: q = 3'b100;
	13'd4988: q = 3'b100;
	13'd4989: q = 3'b100;
	13'd4990: q = 3'b100;
	13'd4991: q = 3'b100;
	13'd4992: q = 3'b100;
	13'd4993: q = 3'b100;
	13'd4994: q = 3'b100;
	13'd4995: q = 3'b100;
	13'd4996: q = 3'b100;
	13'd4997: q = 3'b100;
	13'd4998: q = 3'b100;
	13'd4999: q = 3'b100;
	13'd5000: q = 3'b100;
	13'd5001: q = 3'b100;
	13'd5002: q = 3'b100;
	13'd5003: q = 3'b100;
	13'd5004: q = 3'b100;
	13'd5005: q = 3'b100;
	13'd5006: q = 3'b100;
	13'd5007: q = 3'b100;
	13'd5008: q = 3'b100;
	13'd5009: q = 3'b100;
	13'd5010: q = 3'b000;
	13'd5011: q = 3'b000;
	13'd5012: q = 3'b111;
	13'd5013: q = 3'b111;
	13'd5014: q = 3'b100;
	13'd5015: q = 3'b100;
	13'd5016: q = 3'b100;
	13'd5017: q = 3'b100;
	13'd5018: q = 3'b100;
	13'd5019: q = 3'b100;
	13'd5020: q = 3'b100;
	13'd5021: q = 3'b100;
	13'd5022: q = 3'b100;
	13'd5023: q = 3'b100;
	13'd5024: q = 3'b100;
	13'd5025: q = 3'b100;
	13'd5026: q = 3'b100;
	13'd5027: q = 3'b100;
	13'd5028: q = 3'b100;
	13'd5029: q = 3'b100;
	13'd5030: q = 3'b100;
	13'd5031: q = 3'b100;
	13'd5032: q = 3'b100;
	13'd5033: q = 3'b100;
	13'd5034: q = 3'b100;
	13'd5035: q = 3'b100;
	13'd5036: q = 3'b100;
	13'd5037: q = 3'b100;
	13'd5038: q = 3'b100;
	13'd5039: q = 3'b100;
	13'd5040: q = 3'b100;
	13'd5041: q = 3'b100;
	13'd5042: q = 3'b000;
	13'd5043: q = 3'b000;
	13'd5044: q = 3'b111;
	13'd5045: q = 3'b111;
	13'd5046: q = 3'b100;
	13'd5047: q = 3'b100;
	13'd5048: q = 3'b100;
	13'd5049: q = 3'b100;
	13'd5050: q = 3'b100;
	13'd5051: q = 3'b100;
	13'd5052: q = 3'b100;
	13'd5053: q = 3'b100;
	13'd5054: q = 3'b100;
	13'd5055: q = 3'b100;
	13'd5056: q = 3'b000;
	13'd5057: q = 3'b000;
	13'd5058: q = 3'b000;
	13'd5059: q = 3'b000;
	13'd5060: q = 3'b000;
	13'd5061: q = 3'b000;
	13'd5062: q = 3'b000;
	13'd5063: q = 3'b000;
	13'd5064: q = 3'b000;
	13'd5065: q = 3'b000;
	13'd5066: q = 3'b000;
	13'd5067: q = 3'b000;
	13'd5068: q = 3'b000;
	13'd5069: q = 3'b000;
	13'd5070: q = 3'b000;
	13'd5071: q = 3'b000;
	13'd5072: q = 3'b000;
	13'd5073: q = 3'b000;
	13'd5074: q = 3'b000;
	13'd5075: q = 3'b000;
	13'd5076: q = 3'b000;
	13'd5077: q = 3'b000;
	13'd5078: q = 3'b000;
	13'd5079: q = 3'b000;
	13'd5080: q = 3'b000;
	13'd5081: q = 3'b000;
	13'd5082: q = 3'b000;
	13'd5083: q = 3'b000;
	13'd5084: q = 3'b000;
	13'd5085: q = 3'b000;
	13'd5086: q = 3'b000;
	13'd5087: q = 3'b000;
	13'd5088: q = 3'b000;
	13'd5089: q = 3'b000;
	13'd5090: q = 3'b000;
	13'd5091: q = 3'b000;
	13'd5092: q = 3'b000;
	13'd5093: q = 3'b000;
	13'd5094: q = 3'b000;
	13'd5095: q = 3'b000;
	13'd5096: q = 3'b000;
	13'd5097: q = 3'b000;
	13'd5098: q = 3'b000;
	13'd5099: q = 3'b000;
	13'd5100: q = 3'b000;
	13'd5101: q = 3'b000;
	13'd5102: q = 3'b000;
	13'd5103: q = 3'b000;
	13'd5104: q = 3'b000;
	13'd5105: q = 3'b000;
	13'd5106: q = 3'b000;
	13'd5107: q = 3'b000;
	13'd5108: q = 3'b000;
	13'd5109: q = 3'b000;
	13'd5110: q = 3'b000;
	13'd5111: q = 3'b000;
	13'd5112: q = 3'b000;
	13'd5113: q = 3'b000;
	13'd5114: q = 3'b000;
	13'd5115: q = 3'b000;
	13'd5116: q = 3'b000;
	13'd5117: q = 3'b000;
	13'd5118: q = 3'b000;
	13'd5119: q = 3'b000;
	13'd5120: q = 3'b000;
	13'd5121: q = 3'b000;
	13'd5122: q = 3'b000;
	13'd5123: q = 3'b000;
	13'd5124: q = 3'b000;
	13'd5125: q = 3'b000;
	13'd5126: q = 3'b000;
	13'd5127: q = 3'b000;
	13'd5128: q = 3'b000;
	13'd5129: q = 3'b000;
	13'd5130: q = 3'b111;
	13'd5131: q = 3'b111;
	13'd5132: q = 3'b111;
	13'd5133: q = 3'b111;
	13'd5134: q = 3'b111;
	13'd5135: q = 3'b111;
	13'd5136: q = 3'b111;
	13'd5137: q = 3'b111;
	13'd5138: q = 3'b111;
	13'd5139: q = 3'b111;
	13'd5140: q = 3'b111;
	13'd5141: q = 3'b111;
	13'd5142: q = 3'b000;
	13'd5143: q = 3'b000;
	13'd5144: q = 3'b000;
	13'd5145: q = 3'b000;
	13'd5146: q = 3'b000;
	13'd5147: q = 3'b000;
	13'd5148: q = 3'b000;
	13'd5149: q = 3'b000;
	13'd5150: q = 3'b000;
	13'd5151: q = 3'b000;
	13'd5152: q = 3'b000;
	13'd5153: q = 3'b000;
	13'd5154: q = 3'b000;
	13'd5155: q = 3'b000;
	13'd5156: q = 3'b000;
	13'd5157: q = 3'b000;
	13'd5158: q = 3'b000;
	13'd5159: q = 3'b000;
	13'd5160: q = 3'b000;
	13'd5161: q = 3'b000;
	13'd5162: q = 3'b111;
	13'd5163: q = 3'b111;
	13'd5164: q = 3'b111;
	13'd5165: q = 3'b111;
	13'd5166: q = 3'b111;
	13'd5167: q = 3'b111;
	13'd5168: q = 3'b111;
	13'd5169: q = 3'b111;
	13'd5170: q = 3'b111;
	13'd5171: q = 3'b111;
	13'd5172: q = 3'b111;
	13'd5173: q = 3'b111;
	13'd5174: q = 3'b000;
	13'd5175: q = 3'b000;
	13'd5176: q = 3'b000;
	13'd5177: q = 3'b000;
	13'd5178: q = 3'b000;
	13'd5179: q = 3'b000;
	13'd5180: q = 3'b000;
	13'd5181: q = 3'b000;
	13'd5182: q = 3'b000;
	13'd5183: q = 3'b000;
	13'd5184: q = 3'b000;
	13'd5185: q = 3'b000;
	13'd5186: q = 3'b000;
	13'd5187: q = 3'b000;
	13'd5188: q = 3'b000;
	13'd5189: q = 3'b000;
	13'd5190: q = 3'b000;
	13'd5191: q = 3'b000;
	13'd5192: q = 3'b111;
	13'd5193: q = 3'b111;
	13'd5194: q = 3'b111;
	13'd5195: q = 3'b111;
	13'd5196: q = 3'b111;
	13'd5197: q = 3'b111;
	13'd5198: q = 3'b111;
	13'd5199: q = 3'b111;
	13'd5200: q = 3'b111;
	13'd5201: q = 3'b111;
	13'd5202: q = 3'b111;
	13'd5203: q = 3'b111;
	13'd5204: q = 3'b111;
	13'd5205: q = 3'b111;
	13'd5206: q = 3'b111;
	13'd5207: q = 3'b111;
	13'd5208: q = 3'b000;
	13'd5209: q = 3'b000;
	13'd5210: q = 3'b000;
	13'd5211: q = 3'b000;
	13'd5212: q = 3'b000;
	13'd5213: q = 3'b000;
	13'd5214: q = 3'b000;
	13'd5215: q = 3'b000;
	13'd5216: q = 3'b000;
	13'd5217: q = 3'b000;
	13'd5218: q = 3'b000;
	13'd5219: q = 3'b000;
	13'd5220: q = 3'b000;
	13'd5221: q = 3'b000;
	13'd5222: q = 3'b000;
	13'd5223: q = 3'b000;
	13'd5224: q = 3'b111;
	13'd5225: q = 3'b111;
	13'd5226: q = 3'b111;
	13'd5227: q = 3'b111;
	13'd5228: q = 3'b111;
	13'd5229: q = 3'b111;
	13'd5230: q = 3'b111;
	13'd5231: q = 3'b111;
	13'd5232: q = 3'b111;
	13'd5233: q = 3'b111;
	13'd5234: q = 3'b111;
	13'd5235: q = 3'b111;
	13'd5236: q = 3'b111;
	13'd5237: q = 3'b111;
	13'd5238: q = 3'b111;
	13'd5239: q = 3'b111;
	13'd5240: q = 3'b000;
	13'd5241: q = 3'b000;
	13'd5242: q = 3'b000;
	13'd5243: q = 3'b000;
	13'd5244: q = 3'b000;
	13'd5245: q = 3'b000;
	13'd5246: q = 3'b000;
	13'd5247: q = 3'b000;
	13'd5248: q = 3'b000;
	13'd5249: q = 3'b000;
	13'd5250: q = 3'b000;
	13'd5251: q = 3'b000;
	13'd5252: q = 3'b000;
	13'd5253: q = 3'b000;
	13'd5254: q = 3'b000;
	13'd5255: q = 3'b000;
	13'd5256: q = 3'b111;
	13'd5257: q = 3'b111;
	13'd5258: q = 3'b100;
	13'd5259: q = 3'b100;
	13'd5260: q = 3'b000;
	13'd5261: q = 3'b000;
	13'd5262: q = 3'b100;
	13'd5263: q = 3'b100;
	13'd5264: q = 3'b100;
	13'd5265: q = 3'b100;
	13'd5266: q = 3'b000;
	13'd5267: q = 3'b000;
	13'd5268: q = 3'b100;
	13'd5269: q = 3'b100;
	13'd5270: q = 3'b111;
	13'd5271: q = 3'b111;
	13'd5272: q = 3'b000;
	13'd5273: q = 3'b000;
	13'd5274: q = 3'b000;
	13'd5275: q = 3'b000;
	13'd5276: q = 3'b000;
	13'd5277: q = 3'b000;
	13'd5278: q = 3'b000;
	13'd5279: q = 3'b000;
	13'd5280: q = 3'b000;
	13'd5281: q = 3'b000;
	13'd5282: q = 3'b000;
	13'd5283: q = 3'b000;
	13'd5284: q = 3'b000;
	13'd5285: q = 3'b000;
	13'd5286: q = 3'b000;
	13'd5287: q = 3'b000;
	13'd5288: q = 3'b111;
	13'd5289: q = 3'b111;
	13'd5290: q = 3'b100;
	13'd5291: q = 3'b100;
	13'd5292: q = 3'b000;
	13'd5293: q = 3'b000;
	13'd5294: q = 3'b100;
	13'd5295: q = 3'b100;
	13'd5296: q = 3'b100;
	13'd5297: q = 3'b100;
	13'd5298: q = 3'b000;
	13'd5299: q = 3'b000;
	13'd5300: q = 3'b100;
	13'd5301: q = 3'b100;
	13'd5302: q = 3'b111;
	13'd5303: q = 3'b111;
	13'd5304: q = 3'b000;
	13'd5305: q = 3'b000;
	13'd5306: q = 3'b000;
	13'd5307: q = 3'b000;
	13'd5308: q = 3'b000;
	13'd5309: q = 3'b000;
	13'd5310: q = 3'b000;
	13'd5311: q = 3'b000;
	13'd5312: q = 3'b000;
	13'd5313: q = 3'b000;
	13'd5314: q = 3'b000;
	13'd5315: q = 3'b000;
	13'd5316: q = 3'b000;
	13'd5317: q = 3'b000;
	13'd5318: q = 3'b000;
	13'd5319: q = 3'b000;
	13'd5320: q = 3'b111;
	13'd5321: q = 3'b111;
	13'd5322: q = 3'b100;
	13'd5323: q = 3'b100;
	13'd5324: q = 3'b000;
	13'd5325: q = 3'b000;
	13'd5326: q = 3'b100;
	13'd5327: q = 3'b100;
	13'd5328: q = 3'b100;
	13'd5329: q = 3'b100;
	13'd5330: q = 3'b000;
	13'd5331: q = 3'b000;
	13'd5332: q = 3'b100;
	13'd5333: q = 3'b100;
	13'd5334: q = 3'b111;
	13'd5335: q = 3'b111;
	13'd5336: q = 3'b000;
	13'd5337: q = 3'b000;
	13'd5338: q = 3'b000;
	13'd5339: q = 3'b000;
	13'd5340: q = 3'b000;
	13'd5341: q = 3'b000;
	13'd5342: q = 3'b000;
	13'd5343: q = 3'b000;
	13'd5344: q = 3'b000;
	13'd5345: q = 3'b000;
	13'd5346: q = 3'b000;
	13'd5347: q = 3'b000;
	13'd5348: q = 3'b000;
	13'd5349: q = 3'b000;
	13'd5350: q = 3'b000;
	13'd5351: q = 3'b000;
	13'd5352: q = 3'b111;
	13'd5353: q = 3'b111;
	13'd5354: q = 3'b100;
	13'd5355: q = 3'b100;
	13'd5356: q = 3'b000;
	13'd5357: q = 3'b000;
	13'd5358: q = 3'b100;
	13'd5359: q = 3'b100;
	13'd5360: q = 3'b100;
	13'd5361: q = 3'b100;
	13'd5362: q = 3'b000;
	13'd5363: q = 3'b000;
	13'd5364: q = 3'b100;
	13'd5365: q = 3'b100;
	13'd5366: q = 3'b111;
	13'd5367: q = 3'b111;
	13'd5368: q = 3'b000;
	13'd5369: q = 3'b000;
	13'd5370: q = 3'b000;
	13'd5371: q = 3'b000;
	13'd5372: q = 3'b000;
	13'd5373: q = 3'b000;
	13'd5374: q = 3'b000;
	13'd5375: q = 3'b000;
	13'd5376: q = 3'b000;
	13'd5377: q = 3'b000;
	13'd5378: q = 3'b000;
	13'd5379: q = 3'b000;
	13'd5380: q = 3'b000;
	13'd5381: q = 3'b000;
	13'd5382: q = 3'b000;
	13'd5383: q = 3'b000;
	13'd5384: q = 3'b111;
	13'd5385: q = 3'b111;
	13'd5386: q = 3'b111;
	13'd5387: q = 3'b111;
	13'd5388: q = 3'b111;
	13'd5389: q = 3'b111;
	13'd5390: q = 3'b111;
	13'd5391: q = 3'b111;
	13'd5392: q = 3'b111;
	13'd5393: q = 3'b111;
	13'd5394: q = 3'b111;
	13'd5395: q = 3'b111;
	13'd5396: q = 3'b111;
	13'd5397: q = 3'b111;
	13'd5398: q = 3'b111;
	13'd5399: q = 3'b111;
	13'd5400: q = 3'b000;
	13'd5401: q = 3'b000;
	13'd5402: q = 3'b000;
	13'd5403: q = 3'b000;
	13'd5404: q = 3'b000;
	13'd5405: q = 3'b000;
	13'd5406: q = 3'b000;
	13'd5407: q = 3'b000;
	13'd5408: q = 3'b000;
	13'd5409: q = 3'b000;
	13'd5410: q = 3'b000;
	13'd5411: q = 3'b000;
	13'd5412: q = 3'b000;
	13'd5413: q = 3'b000;
	13'd5414: q = 3'b000;
	13'd5415: q = 3'b000;
	13'd5416: q = 3'b111;
	13'd5417: q = 3'b111;
	13'd5418: q = 3'b111;
	13'd5419: q = 3'b111;
	13'd5420: q = 3'b111;
	13'd5421: q = 3'b111;
	13'd5422: q = 3'b111;
	13'd5423: q = 3'b111;
	13'd5424: q = 3'b111;
	13'd5425: q = 3'b111;
	13'd5426: q = 3'b111;
	13'd5427: q = 3'b111;
	13'd5428: q = 3'b111;
	13'd5429: q = 3'b111;
	13'd5430: q = 3'b111;
	13'd5431: q = 3'b111;
	13'd5432: q = 3'b000;
	13'd5433: q = 3'b000;
	13'd5434: q = 3'b000;
	13'd5435: q = 3'b000;
	13'd5436: q = 3'b000;
	13'd5437: q = 3'b000;
	13'd5438: q = 3'b000;
	13'd5439: q = 3'b000;
	13'd5440: q = 3'b000;
	13'd5441: q = 3'b000;
	13'd5442: q = 3'b000;
	13'd5443: q = 3'b000;
	13'd5444: q = 3'b000;
	13'd5445: q = 3'b000;
	13'd5446: q = 3'b000;
	13'd5447: q = 3'b000;
	13'd5448: q = 3'b000;
	13'd5449: q = 3'b000;
	13'd5450: q = 3'b111;
	13'd5451: q = 3'b111;
	13'd5452: q = 3'b111;
	13'd5453: q = 3'b111;
	13'd5454: q = 3'b111;
	13'd5455: q = 3'b111;
	13'd5456: q = 3'b111;
	13'd5457: q = 3'b111;
	13'd5458: q = 3'b111;
	13'd5459: q = 3'b111;
	13'd5460: q = 3'b111;
	13'd5461: q = 3'b111;
	13'd5462: q = 3'b000;
	13'd5463: q = 3'b000;
	13'd5464: q = 3'b000;
	13'd5465: q = 3'b000;
	13'd5466: q = 3'b000;
	13'd5467: q = 3'b000;
	13'd5468: q = 3'b000;
	13'd5469: q = 3'b000;
	13'd5470: q = 3'b000;
	13'd5471: q = 3'b000;
	13'd5472: q = 3'b000;
	13'd5473: q = 3'b000;
	13'd5474: q = 3'b000;
	13'd5475: q = 3'b000;
	13'd5476: q = 3'b000;
	13'd5477: q = 3'b000;
	13'd5478: q = 3'b000;
	13'd5479: q = 3'b000;
	13'd5480: q = 3'b000;
	13'd5481: q = 3'b000;
	13'd5482: q = 3'b111;
	13'd5483: q = 3'b111;
	13'd5484: q = 3'b111;
	13'd5485: q = 3'b111;
	13'd5486: q = 3'b111;
	13'd5487: q = 3'b111;
	13'd5488: q = 3'b111;
	13'd5489: q = 3'b111;
	13'd5490: q = 3'b111;
	13'd5491: q = 3'b111;
	13'd5492: q = 3'b111;
	13'd5493: q = 3'b111;
	13'd5494: q = 3'b000;
	13'd5495: q = 3'b000;
	13'd5496: q = 3'b000;
	13'd5497: q = 3'b000;
	13'd5498: q = 3'b000;
	13'd5499: q = 3'b000;
	13'd5500: q = 3'b000;
	13'd5501: q = 3'b000;
	13'd5502: q = 3'b000;
	13'd5503: q = 3'b000;
	13'd5504: q = 3'b000;
	13'd5505: q = 3'b000;
	13'd5506: q = 3'b000;
	13'd5507: q = 3'b000;
	13'd5508: q = 3'b000;
	13'd5509: q = 3'b000;
	13'd5510: q = 3'b000;
	13'd5511: q = 3'b000;
	13'd5512: q = 3'b000;
	13'd5513: q = 3'b000;
	13'd5514: q = 3'b000;
	13'd5515: q = 3'b000;
	13'd5516: q = 3'b011;
	13'd5517: q = 3'b011;
	13'd5518: q = 3'b011;
	13'd5519: q = 3'b011;
	13'd5520: q = 3'b011;
	13'd5521: q = 3'b011;
	13'd5522: q = 3'b011;
	13'd5523: q = 3'b011;
	13'd5524: q = 3'b000;
	13'd5525: q = 3'b000;
	13'd5526: q = 3'b000;
	13'd5527: q = 3'b000;
	13'd5528: q = 3'b000;
	13'd5529: q = 3'b000;
	13'd5530: q = 3'b000;
	13'd5531: q = 3'b000;
	13'd5532: q = 3'b000;
	13'd5533: q = 3'b000;
	13'd5534: q = 3'b000;
	13'd5535: q = 3'b000;
	13'd5536: q = 3'b000;
	13'd5537: q = 3'b000;
	13'd5538: q = 3'b000;
	13'd5539: q = 3'b000;
	13'd5540: q = 3'b000;
	13'd5541: q = 3'b000;
	13'd5542: q = 3'b000;
	13'd5543: q = 3'b000;
	13'd5544: q = 3'b000;
	13'd5545: q = 3'b000;
	13'd5546: q = 3'b000;
	13'd5547: q = 3'b000;
	13'd5548: q = 3'b011;
	13'd5549: q = 3'b011;
	13'd5550: q = 3'b011;
	13'd5551: q = 3'b011;
	13'd5552: q = 3'b011;
	13'd5553: q = 3'b011;
	13'd5554: q = 3'b011;
	13'd5555: q = 3'b011;
	13'd5556: q = 3'b000;
	13'd5557: q = 3'b000;
	13'd5558: q = 3'b000;
	13'd5559: q = 3'b000;
	13'd5560: q = 3'b000;
	13'd5561: q = 3'b000;
	13'd5562: q = 3'b000;
	13'd5563: q = 3'b000;
	13'd5564: q = 3'b000;
	13'd5565: q = 3'b000;
	13'd5566: q = 3'b000;
	13'd5567: q = 3'b000;
	13'd5568: q = 3'b000;
	13'd5569: q = 3'b000;
	13'd5570: q = 3'b000;
	13'd5571: q = 3'b000;
	13'd5572: q = 3'b000;
	13'd5573: q = 3'b000;
	13'd5574: q = 3'b000;
	13'd5575: q = 3'b000;
	13'd5576: q = 3'b111;
	13'd5577: q = 3'b111;
	13'd5578: q = 3'b111;
	13'd5579: q = 3'b111;
	13'd5580: q = 3'b011;
	13'd5581: q = 3'b011;
	13'd5582: q = 3'b011;
	13'd5583: q = 3'b011;
	13'd5584: q = 3'b011;
	13'd5585: q = 3'b011;
	13'd5586: q = 3'b011;
	13'd5587: q = 3'b011;
	13'd5588: q = 3'b111;
	13'd5589: q = 3'b111;
	13'd5590: q = 3'b111;
	13'd5591: q = 3'b111;
	13'd5592: q = 3'b000;
	13'd5593: q = 3'b000;
	13'd5594: q = 3'b000;
	13'd5595: q = 3'b000;
	13'd5596: q = 3'b000;
	13'd5597: q = 3'b000;
	13'd5598: q = 3'b000;
	13'd5599: q = 3'b000;
	13'd5600: q = 3'b000;
	13'd5601: q = 3'b000;
	13'd5602: q = 3'b000;
	13'd5603: q = 3'b000;
	13'd5604: q = 3'b000;
	13'd5605: q = 3'b000;
	13'd5606: q = 3'b000;
	13'd5607: q = 3'b000;
	13'd5608: q = 3'b111;
	13'd5609: q = 3'b111;
	13'd5610: q = 3'b111;
	13'd5611: q = 3'b111;
	13'd5612: q = 3'b011;
	13'd5613: q = 3'b011;
	13'd5614: q = 3'b011;
	13'd5615: q = 3'b011;
	13'd5616: q = 3'b011;
	13'd5617: q = 3'b011;
	13'd5618: q = 3'b011;
	13'd5619: q = 3'b011;
	13'd5620: q = 3'b111;
	13'd5621: q = 3'b111;
	13'd5622: q = 3'b111;
	13'd5623: q = 3'b111;
	13'd5624: q = 3'b000;
	13'd5625: q = 3'b000;
	13'd5626: q = 3'b000;
	13'd5627: q = 3'b000;
	13'd5628: q = 3'b000;
	13'd5629: q = 3'b000;
	13'd5630: q = 3'b000;
	13'd5631: q = 3'b000;
	13'd5632: q = 3'b000;
	13'd5633: q = 3'b000;
	13'd5634: q = 3'b000;
	13'd5635: q = 3'b000;
	13'd5636: q = 3'b000;
	13'd5637: q = 3'b000;
	13'd5638: q = 3'b111;
	13'd5639: q = 3'b111;
	13'd5640: q = 3'b111;
	13'd5641: q = 3'b111;
	13'd5642: q = 3'b011;
	13'd5643: q = 3'b011;
	13'd5644: q = 3'b011;
	13'd5645: q = 3'b011;
	13'd5646: q = 3'b011;
	13'd5647: q = 3'b011;
	13'd5648: q = 3'b011;
	13'd5649: q = 3'b011;
	13'd5650: q = 3'b011;
	13'd5651: q = 3'b011;
	13'd5652: q = 3'b011;
	13'd5653: q = 3'b011;
	13'd5654: q = 3'b111;
	13'd5655: q = 3'b111;
	13'd5656: q = 3'b111;
	13'd5657: q = 3'b111;
	13'd5658: q = 3'b000;
	13'd5659: q = 3'b000;
	13'd5660: q = 3'b000;
	13'd5661: q = 3'b000;
	13'd5662: q = 3'b000;
	13'd5663: q = 3'b000;
	13'd5664: q = 3'b000;
	13'd5665: q = 3'b000;
	13'd5666: q = 3'b000;
	13'd5667: q = 3'b000;
	13'd5668: q = 3'b000;
	13'd5669: q = 3'b000;
	13'd5670: q = 3'b111;
	13'd5671: q = 3'b111;
	13'd5672: q = 3'b111;
	13'd5673: q = 3'b111;
	13'd5674: q = 3'b011;
	13'd5675: q = 3'b011;
	13'd5676: q = 3'b011;
	13'd5677: q = 3'b011;
	13'd5678: q = 3'b011;
	13'd5679: q = 3'b011;
	13'd5680: q = 3'b011;
	13'd5681: q = 3'b011;
	13'd5682: q = 3'b011;
	13'd5683: q = 3'b011;
	13'd5684: q = 3'b011;
	13'd5685: q = 3'b011;
	13'd5686: q = 3'b111;
	13'd5687: q = 3'b111;
	13'd5688: q = 3'b111;
	13'd5689: q = 3'b111;
	13'd5690: q = 3'b000;
	13'd5691: q = 3'b000;
	13'd5692: q = 3'b000;
	13'd5693: q = 3'b000;
	13'd5694: q = 3'b000;
	13'd5695: q = 3'b000;
	13'd5696: q = 3'b000;
	13'd5697: q = 3'b000;
	13'd5698: q = 3'b000;
	13'd5699: q = 3'b000;
	13'd5700: q = 3'b100;
	13'd5701: q = 3'b100;
	13'd5702: q = 3'b100;
	13'd5703: q = 3'b100;
	13'd5704: q = 3'b111;
	13'd5705: q = 3'b111;
	13'd5706: q = 3'b011;
	13'd5707: q = 3'b011;
	13'd5708: q = 3'b011;
	13'd5709: q = 3'b011;
	13'd5710: q = 3'b011;
	13'd5711: q = 3'b011;
	13'd5712: q = 3'b011;
	13'd5713: q = 3'b011;
	13'd5714: q = 3'b011;
	13'd5715: q = 3'b011;
	13'd5716: q = 3'b011;
	13'd5717: q = 3'b011;
	13'd5718: q = 3'b111;
	13'd5719: q = 3'b111;
	13'd5720: q = 3'b100;
	13'd5721: q = 3'b100;
	13'd5722: q = 3'b100;
	13'd5723: q = 3'b100;
	13'd5724: q = 3'b000;
	13'd5725: q = 3'b000;
	13'd5726: q = 3'b000;
	13'd5727: q = 3'b000;
	13'd5728: q = 3'b000;
	13'd5729: q = 3'b000;
	13'd5730: q = 3'b000;
	13'd5731: q = 3'b000;
	13'd5732: q = 3'b100;
	13'd5733: q = 3'b100;
	13'd5734: q = 3'b100;
	13'd5735: q = 3'b100;
	13'd5736: q = 3'b111;
	13'd5737: q = 3'b111;
	13'd5738: q = 3'b011;
	13'd5739: q = 3'b011;
	13'd5740: q = 3'b011;
	13'd5741: q = 3'b011;
	13'd5742: q = 3'b011;
	13'd5743: q = 3'b011;
	13'd5744: q = 3'b011;
	13'd5745: q = 3'b011;
	13'd5746: q = 3'b011;
	13'd5747: q = 3'b011;
	13'd5748: q = 3'b011;
	13'd5749: q = 3'b011;
	13'd5750: q = 3'b111;
	13'd5751: q = 3'b111;
	13'd5752: q = 3'b100;
	13'd5753: q = 3'b100;
	13'd5754: q = 3'b100;
	13'd5755: q = 3'b100;
	13'd5756: q = 3'b000;
	13'd5757: q = 3'b000;
	13'd5758: q = 3'b000;
	13'd5759: q = 3'b000;
	13'd5760: q = 3'b000;
	13'd5761: q = 3'b000;
	13'd5762: q = 3'b000;
	13'd5763: q = 3'b000;
	13'd5764: q = 3'b100;
	13'd5765: q = 3'b100;
	13'd5766: q = 3'b100;
	13'd5767: q = 3'b100;
	13'd5768: q = 3'b000;
	13'd5769: q = 3'b000;
	13'd5770: q = 3'b011;
	13'd5771: q = 3'b011;
	13'd5772: q = 3'b011;
	13'd5773: q = 3'b011;
	13'd5774: q = 3'b011;
	13'd5775: q = 3'b011;
	13'd5776: q = 3'b011;
	13'd5777: q = 3'b011;
	13'd5778: q = 3'b011;
	13'd5779: q = 3'b011;
	13'd5780: q = 3'b011;
	13'd5781: q = 3'b011;
	13'd5782: q = 3'b000;
	13'd5783: q = 3'b000;
	13'd5784: q = 3'b100;
	13'd5785: q = 3'b100;
	13'd5786: q = 3'b100;
	13'd5787: q = 3'b100;
	13'd5788: q = 3'b000;
	13'd5789: q = 3'b000;
	13'd5790: q = 3'b000;
	13'd5791: q = 3'b000;
	13'd5792: q = 3'b000;
	13'd5793: q = 3'b000;
	13'd5794: q = 3'b000;
	13'd5795: q = 3'b000;
	13'd5796: q = 3'b100;
	13'd5797: q = 3'b100;
	13'd5798: q = 3'b100;
	13'd5799: q = 3'b100;
	13'd5800: q = 3'b000;
	13'd5801: q = 3'b000;
	13'd5802: q = 3'b011;
	13'd5803: q = 3'b011;
	13'd5804: q = 3'b011;
	13'd5805: q = 3'b011;
	13'd5806: q = 3'b011;
	13'd5807: q = 3'b011;
	13'd5808: q = 3'b011;
	13'd5809: q = 3'b011;
	13'd5810: q = 3'b011;
	13'd5811: q = 3'b011;
	13'd5812: q = 3'b011;
	13'd5813: q = 3'b011;
	13'd5814: q = 3'b000;
	13'd5815: q = 3'b000;
	13'd5816: q = 3'b100;
	13'd5817: q = 3'b100;
	13'd5818: q = 3'b100;
	13'd5819: q = 3'b100;
	13'd5820: q = 3'b000;
	13'd5821: q = 3'b000;
	13'd5822: q = 3'b000;
	13'd5823: q = 3'b000;
	13'd5824: q = 3'b000;
	13'd5825: q = 3'b000;
	13'd5826: q = 3'b000;
	13'd5827: q = 3'b000;
	13'd5828: q = 3'b000;
	13'd5829: q = 3'b000;
	13'd5830: q = 3'b000;
	13'd5831: q = 3'b000;
	13'd5832: q = 3'b000;
	13'd5833: q = 3'b000;
	13'd5834: q = 3'b011;
	13'd5835: q = 3'b011;
	13'd5836: q = 3'b011;
	13'd5837: q = 3'b011;
	13'd5838: q = 3'b011;
	13'd5839: q = 3'b011;
	13'd5840: q = 3'b011;
	13'd5841: q = 3'b011;
	13'd5842: q = 3'b011;
	13'd5843: q = 3'b011;
	13'd5844: q = 3'b011;
	13'd5845: q = 3'b011;
	13'd5846: q = 3'b000;
	13'd5847: q = 3'b000;
	13'd5848: q = 3'b000;
	13'd5849: q = 3'b000;
	13'd5850: q = 3'b000;
	13'd5851: q = 3'b000;
	13'd5852: q = 3'b000;
	13'd5853: q = 3'b000;
	13'd5854: q = 3'b000;
	13'd5855: q = 3'b000;
	13'd5856: q = 3'b000;
	13'd5857: q = 3'b000;
	13'd5858: q = 3'b000;
	13'd5859: q = 3'b000;
	13'd5860: q = 3'b000;
	13'd5861: q = 3'b000;
	13'd5862: q = 3'b000;
	13'd5863: q = 3'b000;
	13'd5864: q = 3'b000;
	13'd5865: q = 3'b000;
	13'd5866: q = 3'b011;
	13'd5867: q = 3'b011;
	13'd5868: q = 3'b011;
	13'd5869: q = 3'b011;
	13'd5870: q = 3'b011;
	13'd5871: q = 3'b011;
	13'd5872: q = 3'b011;
	13'd5873: q = 3'b011;
	13'd5874: q = 3'b011;
	13'd5875: q = 3'b011;
	13'd5876: q = 3'b011;
	13'd5877: q = 3'b011;
	13'd5878: q = 3'b000;
	13'd5879: q = 3'b000;
	13'd5880: q = 3'b000;
	13'd5881: q = 3'b000;
	13'd5882: q = 3'b000;
	13'd5883: q = 3'b000;
	13'd5884: q = 3'b000;
	13'd5885: q = 3'b000;
	13'd5886: q = 3'b000;
	13'd5887: q = 3'b000;
	13'd5888: q = 3'b000;
	13'd5889: q = 3'b000;
	13'd5890: q = 3'b000;
	13'd5891: q = 3'b000;
	13'd5892: q = 3'b000;
	13'd5893: q = 3'b000;
	13'd5894: q = 3'b000;
	13'd5895: q = 3'b000;
	13'd5896: q = 3'b000;
	13'd5897: q = 3'b000;
	13'd5898: q = 3'b111;
	13'd5899: q = 3'b111;
	13'd5900: q = 3'b111;
	13'd5901: q = 3'b111;
	13'd5902: q = 3'b011;
	13'd5903: q = 3'b011;
	13'd5904: q = 3'b011;
	13'd5905: q = 3'b011;
	13'd5906: q = 3'b111;
	13'd5907: q = 3'b111;
	13'd5908: q = 3'b111;
	13'd5909: q = 3'b111;
	13'd5910: q = 3'b000;
	13'd5911: q = 3'b000;
	13'd5912: q = 3'b000;
	13'd5913: q = 3'b000;
	13'd5914: q = 3'b000;
	13'd5915: q = 3'b000;
	13'd5916: q = 3'b000;
	13'd5917: q = 3'b000;
	13'd5918: q = 3'b000;
	13'd5919: q = 3'b000;
	13'd5920: q = 3'b000;
	13'd5921: q = 3'b000;
	13'd5922: q = 3'b000;
	13'd5923: q = 3'b000;
	13'd5924: q = 3'b000;
	13'd5925: q = 3'b000;
	13'd5926: q = 3'b000;
	13'd5927: q = 3'b000;
	13'd5928: q = 3'b000;
	13'd5929: q = 3'b000;
	13'd5930: q = 3'b111;
	13'd5931: q = 3'b111;
	13'd5932: q = 3'b111;
	13'd5933: q = 3'b111;
	13'd5934: q = 3'b011;
	13'd5935: q = 3'b011;
	13'd5936: q = 3'b011;
	13'd5937: q = 3'b011;
	13'd5938: q = 3'b111;
	13'd5939: q = 3'b111;
	13'd5940: q = 3'b111;
	13'd5941: q = 3'b111;
	13'd5942: q = 3'b000;
	13'd5943: q = 3'b000;
	13'd5944: q = 3'b000;
	13'd5945: q = 3'b000;
	13'd5946: q = 3'b000;
	13'd5947: q = 3'b000;
	13'd5948: q = 3'b000;
	13'd5949: q = 3'b000;
	13'd5950: q = 3'b000;
	13'd5951: q = 3'b000;
	13'd5952: q = 3'b000;
	13'd5953: q = 3'b000;
	13'd5954: q = 3'b000;
	13'd5955: q = 3'b000;
	13'd5956: q = 3'b000;
	13'd5957: q = 3'b000;
	13'd5958: q = 3'b000;
	13'd5959: q = 3'b000;
	13'd5960: q = 3'b000;
	13'd5961: q = 3'b000;
	13'd5962: q = 3'b111;
	13'd5963: q = 3'b111;
	13'd5964: q = 3'b111;
	13'd5965: q = 3'b111;
	13'd5966: q = 3'b000;
	13'd5967: q = 3'b000;
	13'd5968: q = 3'b000;
	13'd5969: q = 3'b000;
	13'd5970: q = 3'b111;
	13'd5971: q = 3'b111;
	13'd5972: q = 3'b111;
	13'd5973: q = 3'b111;
	13'd5974: q = 3'b000;
	13'd5975: q = 3'b000;
	13'd5976: q = 3'b000;
	13'd5977: q = 3'b000;
	13'd5978: q = 3'b000;
	13'd5979: q = 3'b000;
	13'd5980: q = 3'b000;
	13'd5981: q = 3'b000;
	13'd5982: q = 3'b000;
	13'd5983: q = 3'b000;
	13'd5984: q = 3'b000;
	13'd5985: q = 3'b000;
	13'd5986: q = 3'b000;
	13'd5987: q = 3'b000;
	13'd5988: q = 3'b000;
	13'd5989: q = 3'b000;
	13'd5990: q = 3'b000;
	13'd5991: q = 3'b000;
	13'd5992: q = 3'b000;
	13'd5993: q = 3'b000;
	13'd5994: q = 3'b111;
	13'd5995: q = 3'b111;
	13'd5996: q = 3'b111;
	13'd5997: q = 3'b111;
	13'd5998: q = 3'b000;
	13'd5999: q = 3'b000;
	13'd6000: q = 3'b000;
	13'd6001: q = 3'b000;
	13'd6002: q = 3'b111;
	13'd6003: q = 3'b111;
	13'd6004: q = 3'b111;
	13'd6005: q = 3'b111;
	13'd6006: q = 3'b000;
	13'd6007: q = 3'b000;
	13'd6008: q = 3'b000;
	13'd6009: q = 3'b000;
	13'd6010: q = 3'b000;
	13'd6011: q = 3'b000;
	13'd6012: q = 3'b000;
	13'd6013: q = 3'b000;
	13'd6014: q = 3'b000;
	13'd6015: q = 3'b000;
	13'd6016: q = 3'b000;
	13'd6017: q = 3'b000;
	13'd6018: q = 3'b000;
	13'd6019: q = 3'b000;
	13'd6020: q = 3'b000;
	13'd6021: q = 3'b000;
	13'd6022: q = 3'b000;
	13'd6023: q = 3'b000;
	13'd6024: q = 3'b000;
	13'd6025: q = 3'b000;
	13'd6026: q = 3'b100;
	13'd6027: q = 3'b100;
	13'd6028: q = 3'b100;
	13'd6029: q = 3'b100;
	13'd6030: q = 3'b000;
	13'd6031: q = 3'b000;
	13'd6032: q = 3'b000;
	13'd6033: q = 3'b000;
	13'd6034: q = 3'b100;
	13'd6035: q = 3'b100;
	13'd6036: q = 3'b100;
	13'd6037: q = 3'b100;
	13'd6038: q = 3'b000;
	13'd6039: q = 3'b000;
	13'd6040: q = 3'b000;
	13'd6041: q = 3'b000;
	13'd6042: q = 3'b000;
	13'd6043: q = 3'b000;
	13'd6044: q = 3'b000;
	13'd6045: q = 3'b000;
	13'd6046: q = 3'b000;
	13'd6047: q = 3'b000;
	13'd6048: q = 3'b000;
	13'd6049: q = 3'b000;
	13'd6050: q = 3'b000;
	13'd6051: q = 3'b000;
	13'd6052: q = 3'b000;
	13'd6053: q = 3'b000;
	13'd6054: q = 3'b000;
	13'd6055: q = 3'b000;
	13'd6056: q = 3'b000;
	13'd6057: q = 3'b000;
	13'd6058: q = 3'b100;
	13'd6059: q = 3'b100;
	13'd6060: q = 3'b100;
	13'd6061: q = 3'b100;
	13'd6062: q = 3'b000;
	13'd6063: q = 3'b000;
	13'd6064: q = 3'b000;
	13'd6065: q = 3'b000;
	13'd6066: q = 3'b100;
	13'd6067: q = 3'b100;
	13'd6068: q = 3'b100;
	13'd6069: q = 3'b100;
	13'd6070: q = 3'b000;
	13'd6071: q = 3'b000;
	13'd6072: q = 3'b000;
	13'd6073: q = 3'b000;
	13'd6074: q = 3'b000;
	13'd6075: q = 3'b000;
	13'd6076: q = 3'b000;
	13'd6077: q = 3'b000;
	13'd6078: q = 3'b000;
	13'd6079: q = 3'b000;
	13'd6080: q = 3'b000;
	13'd6081: q = 3'b000;
	13'd6082: q = 3'b000;
	13'd6083: q = 3'b000;
	13'd6084: q = 3'b000;
	13'd6085: q = 3'b000;
	13'd6086: q = 3'b000;
	13'd6087: q = 3'b000;
	13'd6088: q = 3'b000;
	13'd6089: q = 3'b000;
	13'd6090: q = 3'b100;
	13'd6091: q = 3'b100;
	13'd6092: q = 3'b100;
	13'd6093: q = 3'b100;
	13'd6094: q = 3'b000;
	13'd6095: q = 3'b000;
	13'd6096: q = 3'b000;
	13'd6097: q = 3'b000;
	13'd6098: q = 3'b100;
	13'd6099: q = 3'b100;
	13'd6100: q = 3'b100;
	13'd6101: q = 3'b100;
	13'd6102: q = 3'b000;
	13'd6103: q = 3'b000;
	13'd6104: q = 3'b000;
	13'd6105: q = 3'b000;
	13'd6106: q = 3'b000;
	13'd6107: q = 3'b000;
	13'd6108: q = 3'b000;
	13'd6109: q = 3'b000;
	13'd6110: q = 3'b000;
	13'd6111: q = 3'b000;
	13'd6112: q = 3'b000;
	13'd6113: q = 3'b000;
	13'd6114: q = 3'b000;
	13'd6115: q = 3'b000;
	13'd6116: q = 3'b000;
	13'd6117: q = 3'b000;
	13'd6118: q = 3'b000;
	13'd6119: q = 3'b000;
	13'd6120: q = 3'b000;
	13'd6121: q = 3'b000;
	13'd6122: q = 3'b100;
	13'd6123: q = 3'b100;
	13'd6124: q = 3'b100;
	13'd6125: q = 3'b100;
	13'd6126: q = 3'b000;
	13'd6127: q = 3'b000;
	13'd6128: q = 3'b000;
	13'd6129: q = 3'b000;
	13'd6130: q = 3'b100;
	13'd6131: q = 3'b100;
	13'd6132: q = 3'b100;
	13'd6133: q = 3'b100;
	13'd6134: q = 3'b000;
	13'd6135: q = 3'b000;
	13'd6136: q = 3'b000;
	13'd6137: q = 3'b000;
	13'd6138: q = 3'b000;
	13'd6139: q = 3'b000;
	13'd6140: q = 3'b000;
	13'd6141: q = 3'b000;
	13'd6142: q = 3'b000;
	13'd6143: q = 3'b000;
	13'd6144: q = 3'b000;
	13'd6145: q = 3'b000;
	13'd6146: q = 3'b000;
	13'd6147: q = 3'b000;
	13'd6148: q = 3'b000;
	13'd6149: q = 3'b000;
	13'd6150: q = 3'b000;
	13'd6151: q = 3'b000;
	13'd6152: q = 3'b000;
	13'd6153: q = 3'b000;
	13'd6154: q = 3'b000;
	13'd6155: q = 3'b000;
	13'd6156: q = 3'b100;
	13'd6157: q = 3'b100;
	13'd6158: q = 3'b100;
	13'd6159: q = 3'b100;
	13'd6160: q = 3'b100;
	13'd6161: q = 3'b100;
	13'd6162: q = 3'b100;
	13'd6163: q = 3'b100;
	13'd6164: q = 3'b000;
	13'd6165: q = 3'b000;
	13'd6166: q = 3'b000;
	13'd6167: q = 3'b000;
	13'd6168: q = 3'b000;
	13'd6169: q = 3'b000;
	13'd6170: q = 3'b000;
	13'd6171: q = 3'b000;
	13'd6172: q = 3'b000;
	13'd6173: q = 3'b000;
	13'd6174: q = 3'b000;
	13'd6175: q = 3'b000;
	13'd6176: q = 3'b000;
	13'd6177: q = 3'b000;
	13'd6178: q = 3'b000;
	13'd6179: q = 3'b000;
	13'd6180: q = 3'b000;
	13'd6181: q = 3'b000;
	13'd6182: q = 3'b000;
	13'd6183: q = 3'b000;
	13'd6184: q = 3'b000;
	13'd6185: q = 3'b000;
	13'd6186: q = 3'b000;
	13'd6187: q = 3'b000;
	13'd6188: q = 3'b100;
	13'd6189: q = 3'b100;
	13'd6190: q = 3'b100;
	13'd6191: q = 3'b100;
	13'd6192: q = 3'b100;
	13'd6193: q = 3'b100;
	13'd6194: q = 3'b100;
	13'd6195: q = 3'b100;
	13'd6196: q = 3'b000;
	13'd6197: q = 3'b000;
	13'd6198: q = 3'b000;
	13'd6199: q = 3'b000;
	13'd6200: q = 3'b000;
	13'd6201: q = 3'b000;
	13'd6202: q = 3'b000;
	13'd6203: q = 3'b000;
	13'd6204: q = 3'b000;
	13'd6205: q = 3'b000;
	13'd6206: q = 3'b000;
	13'd6207: q = 3'b000;
	13'd6208: q = 3'b000;
	13'd6209: q = 3'b000;
	13'd6210: q = 3'b000;
	13'd6211: q = 3'b000;
	13'd6212: q = 3'b000;
	13'd6213: q = 3'b000;
	13'd6214: q = 3'b000;
	13'd6215: q = 3'b000;
	13'd6216: q = 3'b000;
	13'd6217: q = 3'b000;
	13'd6218: q = 3'b100;
	13'd6219: q = 3'b100;
	13'd6220: q = 3'b100;
	13'd6221: q = 3'b100;
	13'd6222: q = 3'b100;
	13'd6223: q = 3'b100;
	13'd6224: q = 3'b100;
	13'd6225: q = 3'b100;
	13'd6226: q = 3'b100;
	13'd6227: q = 3'b100;
	13'd6228: q = 3'b100;
	13'd6229: q = 3'b100;
	13'd6230: q = 3'b000;
	13'd6231: q = 3'b000;
	13'd6232: q = 3'b000;
	13'd6233: q = 3'b000;
	13'd6234: q = 3'b000;
	13'd6235: q = 3'b000;
	13'd6236: q = 3'b000;
	13'd6237: q = 3'b000;
	13'd6238: q = 3'b000;
	13'd6239: q = 3'b000;
	13'd6240: q = 3'b000;
	13'd6241: q = 3'b000;
	13'd6242: q = 3'b000;
	13'd6243: q = 3'b000;
	13'd6244: q = 3'b000;
	13'd6245: q = 3'b000;
	13'd6246: q = 3'b000;
	13'd6247: q = 3'b000;
	13'd6248: q = 3'b000;
	13'd6249: q = 3'b000;
	13'd6250: q = 3'b100;
	13'd6251: q = 3'b100;
	13'd6252: q = 3'b100;
	13'd6253: q = 3'b100;
	13'd6254: q = 3'b100;
	13'd6255: q = 3'b100;
	13'd6256: q = 3'b100;
	13'd6257: q = 3'b100;
	13'd6258: q = 3'b100;
	13'd6259: q = 3'b100;
	13'd6260: q = 3'b100;
	13'd6261: q = 3'b100;
	13'd6262: q = 3'b000;
	13'd6263: q = 3'b000;
	13'd6264: q = 3'b000;
	13'd6265: q = 3'b000;
	13'd6266: q = 3'b000;
	13'd6267: q = 3'b000;
	13'd6268: q = 3'b000;
	13'd6269: q = 3'b000;
	13'd6270: q = 3'b000;
	13'd6271: q = 3'b000;
	13'd6272: q = 3'b000;
	13'd6273: q = 3'b000;
	13'd6274: q = 3'b000;
	13'd6275: q = 3'b000;
	13'd6276: q = 3'b000;
	13'd6277: q = 3'b000;
	13'd6278: q = 3'b000;
	13'd6279: q = 3'b000;
	13'd6280: q = 3'b100;
	13'd6281: q = 3'b100;
	13'd6282: q = 3'b100;
	13'd6283: q = 3'b100;
	13'd6284: q = 3'b100;
	13'd6285: q = 3'b100;
	13'd6286: q = 3'b100;
	13'd6287: q = 3'b100;
	13'd6288: q = 3'b100;
	13'd6289: q = 3'b100;
	13'd6290: q = 3'b100;
	13'd6291: q = 3'b100;
	13'd6292: q = 3'b100;
	13'd6293: q = 3'b100;
	13'd6294: q = 3'b100;
	13'd6295: q = 3'b100;
	13'd6296: q = 3'b000;
	13'd6297: q = 3'b000;
	13'd6298: q = 3'b000;
	13'd6299: q = 3'b000;
	13'd6300: q = 3'b000;
	13'd6301: q = 3'b000;
	13'd6302: q = 3'b000;
	13'd6303: q = 3'b000;
	13'd6304: q = 3'b000;
	13'd6305: q = 3'b000;
	13'd6306: q = 3'b000;
	13'd6307: q = 3'b000;
	13'd6308: q = 3'b000;
	13'd6309: q = 3'b000;
	13'd6310: q = 3'b000;
	13'd6311: q = 3'b000;
	13'd6312: q = 3'b100;
	13'd6313: q = 3'b100;
	13'd6314: q = 3'b100;
	13'd6315: q = 3'b100;
	13'd6316: q = 3'b100;
	13'd6317: q = 3'b100;
	13'd6318: q = 3'b100;
	13'd6319: q = 3'b100;
	13'd6320: q = 3'b100;
	13'd6321: q = 3'b100;
	13'd6322: q = 3'b100;
	13'd6323: q = 3'b100;
	13'd6324: q = 3'b100;
	13'd6325: q = 3'b100;
	13'd6326: q = 3'b100;
	13'd6327: q = 3'b100;
	13'd6328: q = 3'b000;
	13'd6329: q = 3'b000;
	13'd6330: q = 3'b000;
	13'd6331: q = 3'b000;
	13'd6332: q = 3'b000;
	13'd6333: q = 3'b000;
	13'd6334: q = 3'b000;
	13'd6335: q = 3'b000;
	13'd6336: q = 3'b000;
	13'd6337: q = 3'b000;
	13'd6338: q = 3'b000;
	13'd6339: q = 3'b000;
	13'd6340: q = 3'b000;
	13'd6341: q = 3'b000;
	13'd6342: q = 3'b100;
	13'd6343: q = 3'b100;
	13'd6344: q = 3'b100;
	13'd6345: q = 3'b100;
	13'd6346: q = 3'b100;
	13'd6347: q = 3'b100;
	13'd6348: q = 3'b100;
	13'd6349: q = 3'b100;
	13'd6350: q = 3'b100;
	13'd6351: q = 3'b100;
	13'd6352: q = 3'b100;
	13'd6353: q = 3'b100;
	13'd6354: q = 3'b100;
	13'd6355: q = 3'b100;
	13'd6356: q = 3'b100;
	13'd6357: q = 3'b100;
	13'd6358: q = 3'b100;
	13'd6359: q = 3'b100;
	13'd6360: q = 3'b100;
	13'd6361: q = 3'b100;
	13'd6362: q = 3'b000;
	13'd6363: q = 3'b000;
	13'd6364: q = 3'b000;
	13'd6365: q = 3'b000;
	13'd6366: q = 3'b000;
	13'd6367: q = 3'b000;
	13'd6368: q = 3'b000;
	13'd6369: q = 3'b000;
	13'd6370: q = 3'b000;
	13'd6371: q = 3'b000;
	13'd6372: q = 3'b000;
	13'd6373: q = 3'b000;
	13'd6374: q = 3'b100;
	13'd6375: q = 3'b100;
	13'd6376: q = 3'b100;
	13'd6377: q = 3'b100;
	13'd6378: q = 3'b100;
	13'd6379: q = 3'b100;
	13'd6380: q = 3'b100;
	13'd6381: q = 3'b100;
	13'd6382: q = 3'b100;
	13'd6383: q = 3'b100;
	13'd6384: q = 3'b100;
	13'd6385: q = 3'b100;
	13'd6386: q = 3'b100;
	13'd6387: q = 3'b100;
	13'd6388: q = 3'b100;
	13'd6389: q = 3'b100;
	13'd6390: q = 3'b100;
	13'd6391: q = 3'b100;
	13'd6392: q = 3'b100;
	13'd6393: q = 3'b100;
	13'd6394: q = 3'b000;
	13'd6395: q = 3'b000;
	13'd6396: q = 3'b000;
	13'd6397: q = 3'b000;
	13'd6398: q = 3'b000;
	13'd6399: q = 3'b000;
	13'd6400: q = 3'b000;
	13'd6401: q = 3'b000;
	13'd6402: q = 3'b000;
	13'd6403: q = 3'b000;
	13'd6404: q = 3'b100;
	13'd6405: q = 3'b100;
	13'd6406: q = 3'b111;
	13'd6407: q = 3'b111;
	13'd6408: q = 3'b111;
	13'd6409: q = 3'b111;
	13'd6410: q = 3'b100;
	13'd6411: q = 3'b100;
	13'd6412: q = 3'b100;
	13'd6413: q = 3'b100;
	13'd6414: q = 3'b100;
	13'd6415: q = 3'b100;
	13'd6416: q = 3'b100;
	13'd6417: q = 3'b100;
	13'd6418: q = 3'b100;
	13'd6419: q = 3'b100;
	13'd6420: q = 3'b100;
	13'd6421: q = 3'b100;
	13'd6422: q = 3'b111;
	13'd6423: q = 3'b111;
	13'd6424: q = 3'b111;
	13'd6425: q = 3'b111;
	13'd6426: q = 3'b100;
	13'd6427: q = 3'b100;
	13'd6428: q = 3'b000;
	13'd6429: q = 3'b000;
	13'd6430: q = 3'b000;
	13'd6431: q = 3'b000;
	13'd6432: q = 3'b000;
	13'd6433: q = 3'b000;
	13'd6434: q = 3'b000;
	13'd6435: q = 3'b000;
	13'd6436: q = 3'b100;
	13'd6437: q = 3'b100;
	13'd6438: q = 3'b111;
	13'd6439: q = 3'b111;
	13'd6440: q = 3'b111;
	13'd6441: q = 3'b111;
	13'd6442: q = 3'b100;
	13'd6443: q = 3'b100;
	13'd6444: q = 3'b100;
	13'd6445: q = 3'b100;
	13'd6446: q = 3'b100;
	13'd6447: q = 3'b100;
	13'd6448: q = 3'b100;
	13'd6449: q = 3'b100;
	13'd6450: q = 3'b100;
	13'd6451: q = 3'b100;
	13'd6452: q = 3'b100;
	13'd6453: q = 3'b100;
	13'd6454: q = 3'b111;
	13'd6455: q = 3'b111;
	13'd6456: q = 3'b111;
	13'd6457: q = 3'b111;
	13'd6458: q = 3'b100;
	13'd6459: q = 3'b100;
	13'd6460: q = 3'b000;
	13'd6461: q = 3'b000;
	13'd6462: q = 3'b000;
	13'd6463: q = 3'b000;
	13'd6464: q = 3'b000;
	13'd6465: q = 3'b000;
	13'd6466: q = 3'b100;
	13'd6467: q = 3'b100;
	13'd6468: q = 3'b100;
	13'd6469: q = 3'b100;
	13'd6470: q = 3'b100;
	13'd6471: q = 3'b100;
	13'd6472: q = 3'b110;
	13'd6473: q = 3'b110;
	13'd6474: q = 3'b111;
	13'd6475: q = 3'b111;
	13'd6476: q = 3'b100;
	13'd6477: q = 3'b100;
	13'd6478: q = 3'b100;
	13'd6479: q = 3'b100;
	13'd6480: q = 3'b100;
	13'd6481: q = 3'b100;
	13'd6482: q = 3'b100;
	13'd6483: q = 3'b100;
	13'd6484: q = 3'b111;
	13'd6485: q = 3'b111;
	13'd6486: q = 3'b110;
	13'd6487: q = 3'b110;
	13'd6488: q = 3'b100;
	13'd6489: q = 3'b100;
	13'd6490: q = 3'b100;
	13'd6491: q = 3'b100;
	13'd6492: q = 3'b100;
	13'd6493: q = 3'b100;
	13'd6494: q = 3'b000;
	13'd6495: q = 3'b000;
	13'd6496: q = 3'b000;
	13'd6497: q = 3'b000;
	13'd6498: q = 3'b100;
	13'd6499: q = 3'b100;
	13'd6500: q = 3'b100;
	13'd6501: q = 3'b100;
	13'd6502: q = 3'b100;
	13'd6503: q = 3'b100;
	13'd6504: q = 3'b110;
	13'd6505: q = 3'b110;
	13'd6506: q = 3'b111;
	13'd6507: q = 3'b111;
	13'd6508: q = 3'b100;
	13'd6509: q = 3'b100;
	13'd6510: q = 3'b100;
	13'd6511: q = 3'b100;
	13'd6512: q = 3'b100;
	13'd6513: q = 3'b100;
	13'd6514: q = 3'b100;
	13'd6515: q = 3'b100;
	13'd6516: q = 3'b111;
	13'd6517: q = 3'b111;
	13'd6518: q = 3'b110;
	13'd6519: q = 3'b110;
	13'd6520: q = 3'b100;
	13'd6521: q = 3'b100;
	13'd6522: q = 3'b100;
	13'd6523: q = 3'b100;
	13'd6524: q = 3'b100;
	13'd6525: q = 3'b100;
	13'd6526: q = 3'b000;
	13'd6527: q = 3'b000;
	13'd6528: q = 3'b000;
	13'd6529: q = 3'b000;
	13'd6530: q = 3'b100;
	13'd6531: q = 3'b100;
	13'd6532: q = 3'b100;
	13'd6533: q = 3'b100;
	13'd6534: q = 3'b100;
	13'd6535: q = 3'b100;
	13'd6536: q = 3'b110;
	13'd6537: q = 3'b110;
	13'd6538: q = 3'b011;
	13'd6539: q = 3'b011;
	13'd6540: q = 3'b111;
	13'd6541: q = 3'b111;
	13'd6542: q = 3'b111;
	13'd6543: q = 3'b111;
	13'd6544: q = 3'b111;
	13'd6545: q = 3'b111;
	13'd6546: q = 3'b111;
	13'd6547: q = 3'b111;
	13'd6548: q = 3'b011;
	13'd6549: q = 3'b011;
	13'd6550: q = 3'b110;
	13'd6551: q = 3'b110;
	13'd6552: q = 3'b100;
	13'd6553: q = 3'b100;
	13'd6554: q = 3'b100;
	13'd6555: q = 3'b100;
	13'd6556: q = 3'b100;
	13'd6557: q = 3'b100;
	13'd6558: q = 3'b000;
	13'd6559: q = 3'b000;
	13'd6560: q = 3'b000;
	13'd6561: q = 3'b000;
	13'd6562: q = 3'b100;
	13'd6563: q = 3'b100;
	13'd6564: q = 3'b100;
	13'd6565: q = 3'b100;
	13'd6566: q = 3'b100;
	13'd6567: q = 3'b100;
	13'd6568: q = 3'b110;
	13'd6569: q = 3'b110;
	13'd6570: q = 3'b011;
	13'd6571: q = 3'b011;
	13'd6572: q = 3'b111;
	13'd6573: q = 3'b111;
	13'd6574: q = 3'b111;
	13'd6575: q = 3'b111;
	13'd6576: q = 3'b111;
	13'd6577: q = 3'b111;
	13'd6578: q = 3'b111;
	13'd6579: q = 3'b111;
	13'd6580: q = 3'b011;
	13'd6581: q = 3'b011;
	13'd6582: q = 3'b110;
	13'd6583: q = 3'b110;
	13'd6584: q = 3'b100;
	13'd6585: q = 3'b100;
	13'd6586: q = 3'b100;
	13'd6587: q = 3'b100;
	13'd6588: q = 3'b100;
	13'd6589: q = 3'b100;
	13'd6590: q = 3'b000;
	13'd6591: q = 3'b000;
	13'd6592: q = 3'b100;
	13'd6593: q = 3'b100;
	13'd6594: q = 3'b100;
	13'd6595: q = 3'b100;
	13'd6596: q = 3'b100;
	13'd6597: q = 3'b100;
	13'd6598: q = 3'b100;
	13'd6599: q = 3'b100;
	13'd6600: q = 3'b110;
	13'd6601: q = 3'b110;
	13'd6602: q = 3'b111;
	13'd6603: q = 3'b111;
	13'd6604: q = 3'b110;
	13'd6605: q = 3'b110;
	13'd6606: q = 3'b100;
	13'd6607: q = 3'b100;
	13'd6608: q = 3'b100;
	13'd6609: q = 3'b100;
	13'd6610: q = 3'b110;
	13'd6611: q = 3'b110;
	13'd6612: q = 3'b111;
	13'd6613: q = 3'b111;
	13'd6614: q = 3'b110;
	13'd6615: q = 3'b110;
	13'd6616: q = 3'b100;
	13'd6617: q = 3'b100;
	13'd6618: q = 3'b100;
	13'd6619: q = 3'b100;
	13'd6620: q = 3'b100;
	13'd6621: q = 3'b100;
	13'd6622: q = 3'b100;
	13'd6623: q = 3'b100;
	13'd6624: q = 3'b100;
	13'd6625: q = 3'b100;
	13'd6626: q = 3'b100;
	13'd6627: q = 3'b100;
	13'd6628: q = 3'b100;
	13'd6629: q = 3'b100;
	13'd6630: q = 3'b100;
	13'd6631: q = 3'b100;
	13'd6632: q = 3'b110;
	13'd6633: q = 3'b110;
	13'd6634: q = 3'b111;
	13'd6635: q = 3'b111;
	13'd6636: q = 3'b110;
	13'd6637: q = 3'b110;
	13'd6638: q = 3'b100;
	13'd6639: q = 3'b100;
	13'd6640: q = 3'b100;
	13'd6641: q = 3'b100;
	13'd6642: q = 3'b110;
	13'd6643: q = 3'b110;
	13'd6644: q = 3'b111;
	13'd6645: q = 3'b111;
	13'd6646: q = 3'b110;
	13'd6647: q = 3'b110;
	13'd6648: q = 3'b100;
	13'd6649: q = 3'b100;
	13'd6650: q = 3'b100;
	13'd6651: q = 3'b100;
	13'd6652: q = 3'b100;
	13'd6653: q = 3'b100;
	13'd6654: q = 3'b100;
	13'd6655: q = 3'b100;
	13'd6656: q = 3'b100;
	13'd6657: q = 3'b100;
	13'd6658: q = 3'b100;
	13'd6659: q = 3'b100;
	13'd6660: q = 3'b100;
	13'd6661: q = 3'b100;
	13'd6662: q = 3'b100;
	13'd6663: q = 3'b100;
	13'd6664: q = 3'b110;
	13'd6665: q = 3'b110;
	13'd6666: q = 3'b110;
	13'd6667: q = 3'b110;
	13'd6668: q = 3'b110;
	13'd6669: q = 3'b110;
	13'd6670: q = 3'b100;
	13'd6671: q = 3'b100;
	13'd6672: q = 3'b100;
	13'd6673: q = 3'b100;
	13'd6674: q = 3'b110;
	13'd6675: q = 3'b110;
	13'd6676: q = 3'b110;
	13'd6677: q = 3'b110;
	13'd6678: q = 3'b110;
	13'd6679: q = 3'b110;
	13'd6680: q = 3'b100;
	13'd6681: q = 3'b100;
	13'd6682: q = 3'b100;
	13'd6683: q = 3'b100;
	13'd6684: q = 3'b100;
	13'd6685: q = 3'b100;
	13'd6686: q = 3'b100;
	13'd6687: q = 3'b100;
	13'd6688: q = 3'b100;
	13'd6689: q = 3'b100;
	13'd6690: q = 3'b100;
	13'd6691: q = 3'b100;
	13'd6692: q = 3'b100;
	13'd6693: q = 3'b100;
	13'd6694: q = 3'b100;
	13'd6695: q = 3'b100;
	13'd6696: q = 3'b110;
	13'd6697: q = 3'b110;
	13'd6698: q = 3'b110;
	13'd6699: q = 3'b110;
	13'd6700: q = 3'b110;
	13'd6701: q = 3'b110;
	13'd6702: q = 3'b100;
	13'd6703: q = 3'b100;
	13'd6704: q = 3'b100;
	13'd6705: q = 3'b100;
	13'd6706: q = 3'b110;
	13'd6707: q = 3'b110;
	13'd6708: q = 3'b110;
	13'd6709: q = 3'b110;
	13'd6710: q = 3'b110;
	13'd6711: q = 3'b110;
	13'd6712: q = 3'b100;
	13'd6713: q = 3'b100;
	13'd6714: q = 3'b100;
	13'd6715: q = 3'b100;
	13'd6716: q = 3'b100;
	13'd6717: q = 3'b100;
	13'd6718: q = 3'b100;
	13'd6719: q = 3'b100;
	13'd6720: q = 3'b100;
	13'd6721: q = 3'b100;
	13'd6722: q = 3'b100;
	13'd6723: q = 3'b100;
	13'd6724: q = 3'b100;
	13'd6725: q = 3'b100;
	13'd6726: q = 3'b100;
	13'd6727: q = 3'b100;
	13'd6728: q = 3'b100;
	13'd6729: q = 3'b100;
	13'd6730: q = 3'b100;
	13'd6731: q = 3'b100;
	13'd6732: q = 3'b100;
	13'd6733: q = 3'b100;
	13'd6734: q = 3'b100;
	13'd6735: q = 3'b100;
	13'd6736: q = 3'b100;
	13'd6737: q = 3'b100;
	13'd6738: q = 3'b100;
	13'd6739: q = 3'b100;
	13'd6740: q = 3'b100;
	13'd6741: q = 3'b100;
	13'd6742: q = 3'b100;
	13'd6743: q = 3'b100;
	13'd6744: q = 3'b100;
	13'd6745: q = 3'b100;
	13'd6746: q = 3'b100;
	13'd6747: q = 3'b100;
	13'd6748: q = 3'b100;
	13'd6749: q = 3'b100;
	13'd6750: q = 3'b100;
	13'd6751: q = 3'b100;
	13'd6752: q = 3'b100;
	13'd6753: q = 3'b100;
	13'd6754: q = 3'b100;
	13'd6755: q = 3'b100;
	13'd6756: q = 3'b100;
	13'd6757: q = 3'b100;
	13'd6758: q = 3'b100;
	13'd6759: q = 3'b100;
	13'd6760: q = 3'b100;
	13'd6761: q = 3'b100;
	13'd6762: q = 3'b100;
	13'd6763: q = 3'b100;
	13'd6764: q = 3'b100;
	13'd6765: q = 3'b100;
	13'd6766: q = 3'b100;
	13'd6767: q = 3'b100;
	13'd6768: q = 3'b100;
	13'd6769: q = 3'b100;
	13'd6770: q = 3'b100;
	13'd6771: q = 3'b100;
	13'd6772: q = 3'b100;
	13'd6773: q = 3'b100;
	13'd6774: q = 3'b100;
	13'd6775: q = 3'b100;
	13'd6776: q = 3'b100;
	13'd6777: q = 3'b100;
	13'd6778: q = 3'b100;
	13'd6779: q = 3'b100;
	13'd6780: q = 3'b100;
	13'd6781: q = 3'b100;
	13'd6782: q = 3'b100;
	13'd6783: q = 3'b100;
	13'd6784: q = 3'b000;
	13'd6785: q = 3'b000;
	13'd6786: q = 3'b100;
	13'd6787: q = 3'b100;
	13'd6788: q = 3'b100;
	13'd6789: q = 3'b100;
	13'd6790: q = 3'b100;
	13'd6791: q = 3'b100;
	13'd6792: q = 3'b100;
	13'd6793: q = 3'b100;
	13'd6794: q = 3'b110;
	13'd6795: q = 3'b110;
	13'd6796: q = 3'b110;
	13'd6797: q = 3'b110;
	13'd6798: q = 3'b110;
	13'd6799: q = 3'b110;
	13'd6800: q = 3'b110;
	13'd6801: q = 3'b110;
	13'd6802: q = 3'b110;
	13'd6803: q = 3'b110;
	13'd6804: q = 3'b110;
	13'd6805: q = 3'b110;
	13'd6806: q = 3'b100;
	13'd6807: q = 3'b100;
	13'd6808: q = 3'b100;
	13'd6809: q = 3'b100;
	13'd6810: q = 3'b100;
	13'd6811: q = 3'b100;
	13'd6812: q = 3'b100;
	13'd6813: q = 3'b100;
	13'd6814: q = 3'b000;
	13'd6815: q = 3'b000;
	13'd6816: q = 3'b000;
	13'd6817: q = 3'b000;
	13'd6818: q = 3'b100;
	13'd6819: q = 3'b100;
	13'd6820: q = 3'b100;
	13'd6821: q = 3'b100;
	13'd6822: q = 3'b100;
	13'd6823: q = 3'b100;
	13'd6824: q = 3'b100;
	13'd6825: q = 3'b100;
	13'd6826: q = 3'b110;
	13'd6827: q = 3'b110;
	13'd6828: q = 3'b110;
	13'd6829: q = 3'b110;
	13'd6830: q = 3'b110;
	13'd6831: q = 3'b110;
	13'd6832: q = 3'b110;
	13'd6833: q = 3'b110;
	13'd6834: q = 3'b110;
	13'd6835: q = 3'b110;
	13'd6836: q = 3'b110;
	13'd6837: q = 3'b110;
	13'd6838: q = 3'b100;
	13'd6839: q = 3'b100;
	13'd6840: q = 3'b100;
	13'd6841: q = 3'b100;
	13'd6842: q = 3'b100;
	13'd6843: q = 3'b100;
	13'd6844: q = 3'b100;
	13'd6845: q = 3'b100;
	13'd6846: q = 3'b000;
	13'd6847: q = 3'b000;
	13'd6848: q = 3'b000;
	13'd6849: q = 3'b000;
	13'd6850: q = 3'b000;
	13'd6851: q = 3'b000;
	13'd6852: q = 3'b000;
	13'd6853: q = 3'b000;
	13'd6854: q = 3'b000;
	13'd6855: q = 3'b000;
	13'd6856: q = 3'b110;
	13'd6857: q = 3'b110;
	13'd6858: q = 3'b110;
	13'd6859: q = 3'b110;
	13'd6860: q = 3'b110;
	13'd6861: q = 3'b110;
	13'd6862: q = 3'b110;
	13'd6863: q = 3'b110;
	13'd6864: q = 3'b110;
	13'd6865: q = 3'b110;
	13'd6866: q = 3'b110;
	13'd6867: q = 3'b110;
	13'd6868: q = 3'b110;
	13'd6869: q = 3'b110;
	13'd6870: q = 3'b110;
	13'd6871: q = 3'b110;
	13'd6872: q = 3'b000;
	13'd6873: q = 3'b000;
	13'd6874: q = 3'b000;
	13'd6875: q = 3'b000;
	13'd6876: q = 3'b000;
	13'd6877: q = 3'b000;
	13'd6878: q = 3'b000;
	13'd6879: q = 3'b000;
	13'd6880: q = 3'b000;
	13'd6881: q = 3'b000;
	13'd6882: q = 3'b000;
	13'd6883: q = 3'b000;
	13'd6884: q = 3'b000;
	13'd6885: q = 3'b000;
	13'd6886: q = 3'b000;
	13'd6887: q = 3'b000;
	13'd6888: q = 3'b110;
	13'd6889: q = 3'b110;
	13'd6890: q = 3'b110;
	13'd6891: q = 3'b110;
	13'd6892: q = 3'b110;
	13'd6893: q = 3'b110;
	13'd6894: q = 3'b110;
	13'd6895: q = 3'b110;
	13'd6896: q = 3'b110;
	13'd6897: q = 3'b110;
	13'd6898: q = 3'b110;
	13'd6899: q = 3'b110;
	13'd6900: q = 3'b110;
	13'd6901: q = 3'b110;
	13'd6902: q = 3'b110;
	13'd6903: q = 3'b110;
	13'd6904: q = 3'b000;
	13'd6905: q = 3'b000;
	13'd6906: q = 3'b000;
	13'd6907: q = 3'b000;
	13'd6908: q = 3'b000;
	13'd6909: q = 3'b000;
	13'd6910: q = 3'b000;
	13'd6911: q = 3'b000;
	13'd6912: q = 3'b000;
	13'd6913: q = 3'b000;
	13'd6914: q = 3'b000;
	13'd6915: q = 3'b000;
	13'd6916: q = 3'b100;
	13'd6917: q = 3'b100;
	13'd6918: q = 3'b100;
	13'd6919: q = 3'b100;
	13'd6920: q = 3'b110;
	13'd6921: q = 3'b110;
	13'd6922: q = 3'b110;
	13'd6923: q = 3'b110;
	13'd6924: q = 3'b110;
	13'd6925: q = 3'b110;
	13'd6926: q = 3'b110;
	13'd6927: q = 3'b110;
	13'd6928: q = 3'b110;
	13'd6929: q = 3'b110;
	13'd6930: q = 3'b110;
	13'd6931: q = 3'b110;
	13'd6932: q = 3'b110;
	13'd6933: q = 3'b110;
	13'd6934: q = 3'b110;
	13'd6935: q = 3'b110;
	13'd6936: q = 3'b100;
	13'd6937: q = 3'b100;
	13'd6938: q = 3'b100;
	13'd6939: q = 3'b100;
	13'd6940: q = 3'b000;
	13'd6941: q = 3'b000;
	13'd6942: q = 3'b000;
	13'd6943: q = 3'b000;
	13'd6944: q = 3'b000;
	13'd6945: q = 3'b000;
	13'd6946: q = 3'b000;
	13'd6947: q = 3'b000;
	13'd6948: q = 3'b100;
	13'd6949: q = 3'b100;
	13'd6950: q = 3'b100;
	13'd6951: q = 3'b100;
	13'd6952: q = 3'b110;
	13'd6953: q = 3'b110;
	13'd6954: q = 3'b110;
	13'd6955: q = 3'b110;
	13'd6956: q = 3'b110;
	13'd6957: q = 3'b110;
	13'd6958: q = 3'b110;
	13'd6959: q = 3'b110;
	13'd6960: q = 3'b110;
	13'd6961: q = 3'b110;
	13'd6962: q = 3'b110;
	13'd6963: q = 3'b110;
	13'd6964: q = 3'b110;
	13'd6965: q = 3'b110;
	13'd6966: q = 3'b110;
	13'd6967: q = 3'b110;
	13'd6968: q = 3'b100;
	13'd6969: q = 3'b100;
	13'd6970: q = 3'b100;
	13'd6971: q = 3'b100;
	13'd6972: q = 3'b000;
	13'd6973: q = 3'b000;
	13'd6974: q = 3'b000;
	13'd6975: q = 3'b000;
	13'd6976: q = 3'b000;
	13'd6977: q = 3'b000;
	13'd6978: q = 3'b100;
	13'd6979: q = 3'b100;
	13'd6980: q = 3'b100;
	13'd6981: q = 3'b100;
	13'd6982: q = 3'b100;
	13'd6983: q = 3'b100;
	13'd6984: q = 3'b100;
	13'd6985: q = 3'b100;
	13'd6986: q = 3'b100;
	13'd6987: q = 3'b100;
	13'd6988: q = 3'b110;
	13'd6989: q = 3'b110;
	13'd6990: q = 3'b110;
	13'd6991: q = 3'b110;
	13'd6992: q = 3'b110;
	13'd6993: q = 3'b110;
	13'd6994: q = 3'b110;
	13'd6995: q = 3'b110;
	13'd6996: q = 3'b100;
	13'd6997: q = 3'b100;
	13'd6998: q = 3'b100;
	13'd6999: q = 3'b100;
	13'd7000: q = 3'b100;
	13'd7001: q = 3'b100;
	13'd7002: q = 3'b100;
	13'd7003: q = 3'b100;
	13'd7004: q = 3'b100;
	13'd7005: q = 3'b100;
	13'd7006: q = 3'b000;
	13'd7007: q = 3'b000;
	13'd7008: q = 3'b000;
	13'd7009: q = 3'b000;
	13'd7010: q = 3'b100;
	13'd7011: q = 3'b100;
	13'd7012: q = 3'b100;
	13'd7013: q = 3'b100;
	13'd7014: q = 3'b100;
	13'd7015: q = 3'b100;
	13'd7016: q = 3'b100;
	13'd7017: q = 3'b100;
	13'd7018: q = 3'b100;
	13'd7019: q = 3'b100;
	13'd7020: q = 3'b110;
	13'd7021: q = 3'b110;
	13'd7022: q = 3'b110;
	13'd7023: q = 3'b110;
	13'd7024: q = 3'b110;
	13'd7025: q = 3'b110;
	13'd7026: q = 3'b110;
	13'd7027: q = 3'b110;
	13'd7028: q = 3'b100;
	13'd7029: q = 3'b100;
	13'd7030: q = 3'b100;
	13'd7031: q = 3'b100;
	13'd7032: q = 3'b100;
	13'd7033: q = 3'b100;
	13'd7034: q = 3'b100;
	13'd7035: q = 3'b100;
	13'd7036: q = 3'b100;
	13'd7037: q = 3'b100;
	13'd7038: q = 3'b000;
	13'd7039: q = 3'b000;
	13'd7040: q = 3'b000;
	13'd7041: q = 3'b000;
	13'd7042: q = 3'b100;
	13'd7043: q = 3'b100;
	13'd7044: q = 3'b100;
	13'd7045: q = 3'b100;
	13'd7046: q = 3'b100;
	13'd7047: q = 3'b100;
	13'd7048: q = 3'b100;
	13'd7049: q = 3'b100;
	13'd7050: q = 3'b100;
	13'd7051: q = 3'b100;
	13'd7052: q = 3'b100;
	13'd7053: q = 3'b100;
	13'd7054: q = 3'b110;
	13'd7055: q = 3'b110;
	13'd7056: q = 3'b110;
	13'd7057: q = 3'b110;
	13'd7058: q = 3'b100;
	13'd7059: q = 3'b100;
	13'd7060: q = 3'b100;
	13'd7061: q = 3'b100;
	13'd7062: q = 3'b100;
	13'd7063: q = 3'b100;
	13'd7064: q = 3'b100;
	13'd7065: q = 3'b100;
	13'd7066: q = 3'b100;
	13'd7067: q = 3'b100;
	13'd7068: q = 3'b100;
	13'd7069: q = 3'b100;
	13'd7070: q = 3'b000;
	13'd7071: q = 3'b000;
	13'd7072: q = 3'b000;
	13'd7073: q = 3'b000;
	13'd7074: q = 3'b100;
	13'd7075: q = 3'b100;
	13'd7076: q = 3'b100;
	13'd7077: q = 3'b100;
	13'd7078: q = 3'b100;
	13'd7079: q = 3'b100;
	13'd7080: q = 3'b100;
	13'd7081: q = 3'b100;
	13'd7082: q = 3'b100;
	13'd7083: q = 3'b100;
	13'd7084: q = 3'b100;
	13'd7085: q = 3'b100;
	13'd7086: q = 3'b110;
	13'd7087: q = 3'b110;
	13'd7088: q = 3'b110;
	13'd7089: q = 3'b110;
	13'd7090: q = 3'b100;
	13'd7091: q = 3'b100;
	13'd7092: q = 3'b100;
	13'd7093: q = 3'b100;
	13'd7094: q = 3'b100;
	13'd7095: q = 3'b100;
	13'd7096: q = 3'b100;
	13'd7097: q = 3'b100;
	13'd7098: q = 3'b100;
	13'd7099: q = 3'b100;
	13'd7100: q = 3'b100;
	13'd7101: q = 3'b100;
	13'd7102: q = 3'b000;
	13'd7103: q = 3'b000;
	13'd7104: q = 3'b000;
	13'd7105: q = 3'b000;
	13'd7106: q = 3'b000;
	13'd7107: q = 3'b000;
	13'd7108: q = 3'b100;
	13'd7109: q = 3'b100;
	13'd7110: q = 3'b100;
	13'd7111: q = 3'b100;
	13'd7112: q = 3'b100;
	13'd7113: q = 3'b100;
	13'd7114: q = 3'b100;
	13'd7115: q = 3'b100;
	13'd7116: q = 3'b100;
	13'd7117: q = 3'b100;
	13'd7118: q = 3'b110;
	13'd7119: q = 3'b110;
	13'd7120: q = 3'b110;
	13'd7121: q = 3'b110;
	13'd7122: q = 3'b100;
	13'd7123: q = 3'b100;
	13'd7124: q = 3'b100;
	13'd7125: q = 3'b100;
	13'd7126: q = 3'b100;
	13'd7127: q = 3'b100;
	13'd7128: q = 3'b100;
	13'd7129: q = 3'b100;
	13'd7130: q = 3'b100;
	13'd7131: q = 3'b100;
	13'd7132: q = 3'b000;
	13'd7133: q = 3'b000;
	13'd7134: q = 3'b000;
	13'd7135: q = 3'b000;
	13'd7136: q = 3'b000;
	13'd7137: q = 3'b000;
	13'd7138: q = 3'b000;
	13'd7139: q = 3'b000;
	13'd7140: q = 3'b100;
	13'd7141: q = 3'b100;
	13'd7142: q = 3'b100;
	13'd7143: q = 3'b100;
	13'd7144: q = 3'b100;
	13'd7145: q = 3'b100;
	13'd7146: q = 3'b100;
	13'd7147: q = 3'b100;
	13'd7148: q = 3'b100;
	13'd7149: q = 3'b100;
	13'd7150: q = 3'b110;
	13'd7151: q = 3'b110;
	13'd7152: q = 3'b110;
	13'd7153: q = 3'b110;
	13'd7154: q = 3'b100;
	13'd7155: q = 3'b100;
	13'd7156: q = 3'b100;
	13'd7157: q = 3'b100;
	13'd7158: q = 3'b100;
	13'd7159: q = 3'b100;
	13'd7160: q = 3'b100;
	13'd7161: q = 3'b100;
	13'd7162: q = 3'b100;
	13'd7163: q = 3'b100;
	13'd7164: q = 3'b000;
	13'd7165: q = 3'b000;
	13'd7166: q = 3'b000;
	13'd7167: q = 3'b000;
	13'd7168: q = 3'b000;
	13'd7169: q = 3'b000;
	13'd7170: q = 3'b000;
	13'd7171: q = 3'b000;
	13'd7172: q = 3'b000;
	13'd7173: q = 3'b000;
	13'd7174: q = 3'b000;
	13'd7175: q = 3'b000;
	13'd7176: q = 3'b000;
	13'd7177: q = 3'b000;
	13'd7178: q = 3'b000;
	13'd7179: q = 3'b000;
	13'd7180: q = 3'b000;
	13'd7181: q = 3'b000;
	13'd7182: q = 3'b000;
	13'd7183: q = 3'b000;
	13'd7184: q = 3'b000;
	13'd7185: q = 3'b000;
	13'd7186: q = 3'b111;
	13'd7187: q = 3'b111;
	13'd7188: q = 3'b111;
	13'd7189: q = 3'b111;
	13'd7190: q = 3'b111;
	13'd7191: q = 3'b111;
	13'd7192: q = 3'b000;
	13'd7193: q = 3'b000;
	13'd7194: q = 3'b111;
	13'd7195: q = 3'b111;
	13'd7196: q = 3'b000;
	13'd7197: q = 3'b000;
	13'd7198: q = 3'b111;
	13'd7199: q = 3'b111;
	13'd7200: q = 3'b000;
	13'd7201: q = 3'b000;
	13'd7202: q = 3'b000;
	13'd7203: q = 3'b000;
	13'd7204: q = 3'b000;
	13'd7205: q = 3'b000;
	13'd7206: q = 3'b000;
	13'd7207: q = 3'b000;
	13'd7208: q = 3'b000;
	13'd7209: q = 3'b000;
	13'd7210: q = 3'b000;
	13'd7211: q = 3'b000;
	13'd7212: q = 3'b000;
	13'd7213: q = 3'b000;
	13'd7214: q = 3'b000;
	13'd7215: q = 3'b000;
	13'd7216: q = 3'b000;
	13'd7217: q = 3'b000;
	13'd7218: q = 3'b111;
	13'd7219: q = 3'b111;
	13'd7220: q = 3'b111;
	13'd7221: q = 3'b111;
	13'd7222: q = 3'b111;
	13'd7223: q = 3'b111;
	13'd7224: q = 3'b000;
	13'd7225: q = 3'b000;
	13'd7226: q = 3'b111;
	13'd7227: q = 3'b111;
	13'd7228: q = 3'b000;
	13'd7229: q = 3'b000;
	13'd7230: q = 3'b111;
	13'd7231: q = 3'b111;
	13'd7232: q = 3'b000;
	13'd7233: q = 3'b000;
	13'd7234: q = 3'b000;
	13'd7235: q = 3'b000;
	13'd7236: q = 3'b000;
	13'd7237: q = 3'b000;
	13'd7238: q = 3'b000;
	13'd7239: q = 3'b000;
	13'd7240: q = 3'b000;
	13'd7241: q = 3'b000;
	13'd7242: q = 3'b100;
	13'd7243: q = 3'b100;
	13'd7244: q = 3'b100;
	13'd7245: q = 3'b100;
	13'd7246: q = 3'b100;
	13'd7247: q = 3'b100;
	13'd7248: q = 3'b111;
	13'd7249: q = 3'b111;
	13'd7250: q = 3'b111;
	13'd7251: q = 3'b111;
	13'd7252: q = 3'b100;
	13'd7253: q = 3'b100;
	13'd7254: q = 3'b100;
	13'd7255: q = 3'b100;
	13'd7256: q = 3'b000;
	13'd7257: q = 3'b000;
	13'd7258: q = 3'b000;
	13'd7259: q = 3'b000;
	13'd7260: q = 3'b000;
	13'd7261: q = 3'b000;
	13'd7262: q = 3'b000;
	13'd7263: q = 3'b000;
	13'd7264: q = 3'b000;
	13'd7265: q = 3'b000;
	13'd7266: q = 3'b000;
	13'd7267: q = 3'b000;
	13'd7268: q = 3'b000;
	13'd7269: q = 3'b000;
	13'd7270: q = 3'b000;
	13'd7271: q = 3'b000;
	13'd7272: q = 3'b000;
	13'd7273: q = 3'b000;
	13'd7274: q = 3'b100;
	13'd7275: q = 3'b100;
	13'd7276: q = 3'b100;
	13'd7277: q = 3'b100;
	13'd7278: q = 3'b100;
	13'd7279: q = 3'b100;
	13'd7280: q = 3'b111;
	13'd7281: q = 3'b111;
	13'd7282: q = 3'b111;
	13'd7283: q = 3'b111;
	13'd7284: q = 3'b100;
	13'd7285: q = 3'b100;
	13'd7286: q = 3'b100;
	13'd7287: q = 3'b100;
	13'd7288: q = 3'b000;
	13'd7289: q = 3'b000;
	13'd7290: q = 3'b000;
	13'd7291: q = 3'b000;
	13'd7292: q = 3'b000;
	13'd7293: q = 3'b000;
	13'd7294: q = 3'b000;
	13'd7295: q = 3'b000;
	13'd7296: q = 3'b000;
	13'd7297: q = 3'b000;
	13'd7298: q = 3'b000;
	13'd7299: q = 3'b000;
	13'd7300: q = 3'b000;
	13'd7301: q = 3'b000;
	13'd7302: q = 3'b100;
	13'd7303: q = 3'b100;
	13'd7304: q = 3'b100;
	13'd7305: q = 3'b100;
	13'd7306: q = 3'b100;
	13'd7307: q = 3'b100;
	13'd7308: q = 3'b100;
	13'd7309: q = 3'b100;
	13'd7310: q = 3'b100;
	13'd7311: q = 3'b100;
	13'd7312: q = 3'b111;
	13'd7313: q = 3'b111;
	13'd7314: q = 3'b100;
	13'd7315: q = 3'b100;
	13'd7316: q = 3'b100;
	13'd7317: q = 3'b100;
	13'd7318: q = 3'b100;
	13'd7319: q = 3'b100;
	13'd7320: q = 3'b100;
	13'd7321: q = 3'b100;
	13'd7322: q = 3'b000;
	13'd7323: q = 3'b000;
	13'd7324: q = 3'b111;
	13'd7325: q = 3'b111;
	13'd7326: q = 3'b000;
	13'd7327: q = 3'b000;
	13'd7328: q = 3'b000;
	13'd7329: q = 3'b000;
	13'd7330: q = 3'b000;
	13'd7331: q = 3'b000;
	13'd7332: q = 3'b000;
	13'd7333: q = 3'b000;
	13'd7334: q = 3'b100;
	13'd7335: q = 3'b100;
	13'd7336: q = 3'b100;
	13'd7337: q = 3'b100;
	13'd7338: q = 3'b100;
	13'd7339: q = 3'b100;
	13'd7340: q = 3'b100;
	13'd7341: q = 3'b100;
	13'd7342: q = 3'b100;
	13'd7343: q = 3'b100;
	13'd7344: q = 3'b111;
	13'd7345: q = 3'b111;
	13'd7346: q = 3'b100;
	13'd7347: q = 3'b100;
	13'd7348: q = 3'b100;
	13'd7349: q = 3'b100;
	13'd7350: q = 3'b100;
	13'd7351: q = 3'b100;
	13'd7352: q = 3'b100;
	13'd7353: q = 3'b100;
	13'd7354: q = 3'b000;
	13'd7355: q = 3'b000;
	13'd7356: q = 3'b111;
	13'd7357: q = 3'b111;
	13'd7358: q = 3'b000;
	13'd7359: q = 3'b000;
	13'd7360: q = 3'b000;
	13'd7361: q = 3'b000;
	13'd7362: q = 3'b000;
	13'd7363: q = 3'b000;
	13'd7364: q = 3'b100;
	13'd7365: q = 3'b100;
	13'd7366: q = 3'b100;
	13'd7367: q = 3'b100;
	13'd7368: q = 3'b111;
	13'd7369: q = 3'b111;
	13'd7370: q = 3'b111;
	13'd7371: q = 3'b111;
	13'd7372: q = 3'b100;
	13'd7373: q = 3'b100;
	13'd7374: q = 3'b100;
	13'd7375: q = 3'b100;
	13'd7376: q = 3'b111;
	13'd7377: q = 3'b111;
	13'd7378: q = 3'b100;
	13'd7379: q = 3'b100;
	13'd7380: q = 3'b100;
	13'd7381: q = 3'b100;
	13'd7382: q = 3'b100;
	13'd7383: q = 3'b100;
	13'd7384: q = 3'b100;
	13'd7385: q = 3'b100;
	13'd7386: q = 3'b100;
	13'd7387: q = 3'b100;
	13'd7388: q = 3'b000;
	13'd7389: q = 3'b000;
	13'd7390: q = 3'b000;
	13'd7391: q = 3'b000;
	13'd7392: q = 3'b000;
	13'd7393: q = 3'b000;
	13'd7394: q = 3'b000;
	13'd7395: q = 3'b000;
	13'd7396: q = 3'b100;
	13'd7397: q = 3'b100;
	13'd7398: q = 3'b100;
	13'd7399: q = 3'b100;
	13'd7400: q = 3'b111;
	13'd7401: q = 3'b111;
	13'd7402: q = 3'b111;
	13'd7403: q = 3'b111;
	13'd7404: q = 3'b100;
	13'd7405: q = 3'b100;
	13'd7406: q = 3'b100;
	13'd7407: q = 3'b100;
	13'd7408: q = 3'b111;
	13'd7409: q = 3'b111;
	13'd7410: q = 3'b100;
	13'd7411: q = 3'b100;
	13'd7412: q = 3'b100;
	13'd7413: q = 3'b100;
	13'd7414: q = 3'b100;
	13'd7415: q = 3'b100;
	13'd7416: q = 3'b100;
	13'd7417: q = 3'b100;
	13'd7418: q = 3'b100;
	13'd7419: q = 3'b100;
	13'd7420: q = 3'b000;
	13'd7421: q = 3'b000;
	13'd7422: q = 3'b000;
	13'd7423: q = 3'b000;
	13'd7424: q = 3'b000;
	13'd7425: q = 3'b000;
	13'd7426: q = 3'b100;
	13'd7427: q = 3'b100;
	13'd7428: q = 3'b100;
	13'd7429: q = 3'b100;
	13'd7430: q = 3'b111;
	13'd7431: q = 3'b111;
	13'd7432: q = 3'b111;
	13'd7433: q = 3'b111;
	13'd7434: q = 3'b100;
	13'd7435: q = 3'b100;
	13'd7436: q = 3'b100;
	13'd7437: q = 3'b100;
	13'd7438: q = 3'b100;
	13'd7439: q = 3'b100;
	13'd7440: q = 3'b100;
	13'd7441: q = 3'b100;
	13'd7442: q = 3'b100;
	13'd7443: q = 3'b100;
	13'd7444: q = 3'b100;
	13'd7445: q = 3'b100;
	13'd7446: q = 3'b100;
	13'd7447: q = 3'b100;
	13'd7448: q = 3'b100;
	13'd7449: q = 3'b100;
	13'd7450: q = 3'b100;
	13'd7451: q = 3'b100;
	13'd7452: q = 3'b100;
	13'd7453: q = 3'b100;
	13'd7454: q = 3'b000;
	13'd7455: q = 3'b000;
	13'd7456: q = 3'b000;
	13'd7457: q = 3'b000;
	13'd7458: q = 3'b100;
	13'd7459: q = 3'b100;
	13'd7460: q = 3'b100;
	13'd7461: q = 3'b100;
	13'd7462: q = 3'b111;
	13'd7463: q = 3'b111;
	13'd7464: q = 3'b111;
	13'd7465: q = 3'b111;
	13'd7466: q = 3'b100;
	13'd7467: q = 3'b100;
	13'd7468: q = 3'b100;
	13'd7469: q = 3'b100;
	13'd7470: q = 3'b100;
	13'd7471: q = 3'b100;
	13'd7472: q = 3'b100;
	13'd7473: q = 3'b100;
	13'd7474: q = 3'b100;
	13'd7475: q = 3'b100;
	13'd7476: q = 3'b100;
	13'd7477: q = 3'b100;
	13'd7478: q = 3'b100;
	13'd7479: q = 3'b100;
	13'd7480: q = 3'b100;
	13'd7481: q = 3'b100;
	13'd7482: q = 3'b100;
	13'd7483: q = 3'b100;
	13'd7484: q = 3'b100;
	13'd7485: q = 3'b100;
	13'd7486: q = 3'b000;
	13'd7487: q = 3'b000;
	13'd7488: q = 3'b000;
	13'd7489: q = 3'b000;
	13'd7490: q = 3'b100;
	13'd7491: q = 3'b100;
	13'd7492: q = 3'b100;
	13'd7493: q = 3'b100;
	13'd7494: q = 3'b111;
	13'd7495: q = 3'b111;
	13'd7496: q = 3'b111;
	13'd7497: q = 3'b111;
	13'd7498: q = 3'b100;
	13'd7499: q = 3'b100;
	13'd7500: q = 3'b100;
	13'd7501: q = 3'b100;
	13'd7502: q = 3'b100;
	13'd7503: q = 3'b100;
	13'd7504: q = 3'b100;
	13'd7505: q = 3'b100;
	13'd7506: q = 3'b100;
	13'd7507: q = 3'b100;
	13'd7508: q = 3'b100;
	13'd7509: q = 3'b100;
	13'd7510: q = 3'b100;
	13'd7511: q = 3'b100;
	13'd7512: q = 3'b100;
	13'd7513: q = 3'b100;
	13'd7514: q = 3'b100;
	13'd7515: q = 3'b100;
	13'd7516: q = 3'b100;
	13'd7517: q = 3'b100;
	13'd7518: q = 3'b000;
	13'd7519: q = 3'b000;
	13'd7520: q = 3'b000;
	13'd7521: q = 3'b000;
	13'd7522: q = 3'b100;
	13'd7523: q = 3'b100;
	13'd7524: q = 3'b100;
	13'd7525: q = 3'b100;
	13'd7526: q = 3'b111;
	13'd7527: q = 3'b111;
	13'd7528: q = 3'b111;
	13'd7529: q = 3'b111;
	13'd7530: q = 3'b100;
	13'd7531: q = 3'b100;
	13'd7532: q = 3'b100;
	13'd7533: q = 3'b100;
	13'd7534: q = 3'b100;
	13'd7535: q = 3'b100;
	13'd7536: q = 3'b100;
	13'd7537: q = 3'b100;
	13'd7538: q = 3'b100;
	13'd7539: q = 3'b100;
	13'd7540: q = 3'b100;
	13'd7541: q = 3'b100;
	13'd7542: q = 3'b100;
	13'd7543: q = 3'b100;
	13'd7544: q = 3'b100;
	13'd7545: q = 3'b100;
	13'd7546: q = 3'b100;
	13'd7547: q = 3'b100;
	13'd7548: q = 3'b100;
	13'd7549: q = 3'b100;
	13'd7550: q = 3'b000;
	13'd7551: q = 3'b000;
	13'd7552: q = 3'b100;
	13'd7553: q = 3'b100;
	13'd7554: q = 3'b100;
	13'd7555: q = 3'b100;
	13'd7556: q = 3'b111;
	13'd7557: q = 3'b111;
	13'd7558: q = 3'b111;
	13'd7559: q = 3'b111;
	13'd7560: q = 3'b100;
	13'd7561: q = 3'b100;
	13'd7562: q = 3'b100;
	13'd7563: q = 3'b100;
	13'd7564: q = 3'b100;
	13'd7565: q = 3'b100;
	13'd7566: q = 3'b100;
	13'd7567: q = 3'b100;
	13'd7568: q = 3'b100;
	13'd7569: q = 3'b100;
	13'd7570: q = 3'b100;
	13'd7571: q = 3'b100;
	13'd7572: q = 3'b100;
	13'd7573: q = 3'b100;
	13'd7574: q = 3'b100;
	13'd7575: q = 3'b100;
	13'd7576: q = 3'b100;
	13'd7577: q = 3'b100;
	13'd7578: q = 3'b100;
	13'd7579: q = 3'b100;
	13'd7580: q = 3'b100;
	13'd7581: q = 3'b100;
	13'd7582: q = 3'b100;
	13'd7583: q = 3'b100;
	13'd7584: q = 3'b100;
	13'd7585: q = 3'b100;
	13'd7586: q = 3'b100;
	13'd7587: q = 3'b100;
	13'd7588: q = 3'b111;
	13'd7589: q = 3'b111;
	13'd7590: q = 3'b111;
	13'd7591: q = 3'b111;
	13'd7592: q = 3'b100;
	13'd7593: q = 3'b100;
	13'd7594: q = 3'b100;
	13'd7595: q = 3'b100;
	13'd7596: q = 3'b100;
	13'd7597: q = 3'b100;
	13'd7598: q = 3'b100;
	13'd7599: q = 3'b100;
	13'd7600: q = 3'b100;
	13'd7601: q = 3'b100;
	13'd7602: q = 3'b100;
	13'd7603: q = 3'b100;
	13'd7604: q = 3'b100;
	13'd7605: q = 3'b100;
	13'd7606: q = 3'b100;
	13'd7607: q = 3'b100;
	13'd7608: q = 3'b100;
	13'd7609: q = 3'b100;
	13'd7610: q = 3'b100;
	13'd7611: q = 3'b100;
	13'd7612: q = 3'b100;
	13'd7613: q = 3'b100;
	13'd7614: q = 3'b100;
	13'd7615: q = 3'b100;
	13'd7616: q = 3'b100;
	13'd7617: q = 3'b100;
	13'd7618: q = 3'b100;
	13'd7619: q = 3'b100;
	13'd7620: q = 3'b111;
	13'd7621: q = 3'b111;
	13'd7622: q = 3'b111;
	13'd7623: q = 3'b111;
	13'd7624: q = 3'b100;
	13'd7625: q = 3'b100;
	13'd7626: q = 3'b100;
	13'd7627: q = 3'b100;
	13'd7628: q = 3'b100;
	13'd7629: q = 3'b100;
	13'd7630: q = 3'b100;
	13'd7631: q = 3'b100;
	13'd7632: q = 3'b100;
	13'd7633: q = 3'b100;
	13'd7634: q = 3'b100;
	13'd7635: q = 3'b100;
	13'd7636: q = 3'b100;
	13'd7637: q = 3'b100;
	13'd7638: q = 3'b100;
	13'd7639: q = 3'b100;
	13'd7640: q = 3'b100;
	13'd7641: q = 3'b100;
	13'd7642: q = 3'b100;
	13'd7643: q = 3'b100;
	13'd7644: q = 3'b100;
	13'd7645: q = 3'b100;
	13'd7646: q = 3'b100;
	13'd7647: q = 3'b100;
	13'd7648: q = 3'b100;
	13'd7649: q = 3'b100;
	13'd7650: q = 3'b100;
	13'd7651: q = 3'b100;
	13'd7652: q = 3'b111;
	13'd7653: q = 3'b111;
	13'd7654: q = 3'b111;
	13'd7655: q = 3'b111;
	13'd7656: q = 3'b100;
	13'd7657: q = 3'b100;
	13'd7658: q = 3'b100;
	13'd7659: q = 3'b100;
	13'd7660: q = 3'b100;
	13'd7661: q = 3'b100;
	13'd7662: q = 3'b100;
	13'd7663: q = 3'b100;
	13'd7664: q = 3'b100;
	13'd7665: q = 3'b100;
	13'd7666: q = 3'b100;
	13'd7667: q = 3'b100;
	13'd7668: q = 3'b100;
	13'd7669: q = 3'b100;
	13'd7670: q = 3'b100;
	13'd7671: q = 3'b100;
	13'd7672: q = 3'b100;
	13'd7673: q = 3'b100;
	13'd7674: q = 3'b100;
	13'd7675: q = 3'b100;
	13'd7676: q = 3'b100;
	13'd7677: q = 3'b100;
	13'd7678: q = 3'b100;
	13'd7679: q = 3'b100;
	13'd7680: q = 3'b100;
	13'd7681: q = 3'b100;
	13'd7682: q = 3'b100;
	13'd7683: q = 3'b100;
	13'd7684: q = 3'b100;
	13'd7685: q = 3'b100;
	13'd7686: q = 3'b100;
	13'd7687: q = 3'b100;
	13'd7688: q = 3'b100;
	13'd7689: q = 3'b100;
	13'd7690: q = 3'b100;
	13'd7691: q = 3'b100;
	13'd7692: q = 3'b100;
	13'd7693: q = 3'b100;
	13'd7694: q = 3'b100;
	13'd7695: q = 3'b100;
	13'd7696: q = 3'b100;
	13'd7697: q = 3'b100;
	13'd7698: q = 3'b100;
	13'd7699: q = 3'b100;
	13'd7700: q = 3'b100;
	13'd7701: q = 3'b100;
	13'd7702: q = 3'b100;
	13'd7703: q = 3'b100;
	13'd7704: q = 3'b100;
	13'd7705: q = 3'b100;
	13'd7706: q = 3'b100;
	13'd7707: q = 3'b100;
	13'd7708: q = 3'b100;
	13'd7709: q = 3'b100;
	13'd7710: q = 3'b100;
	13'd7711: q = 3'b100;
	13'd7712: q = 3'b100;
	13'd7713: q = 3'b100;
	13'd7714: q = 3'b100;
	13'd7715: q = 3'b100;
	13'd7716: q = 3'b100;
	13'd7717: q = 3'b100;
	13'd7718: q = 3'b100;
	13'd7719: q = 3'b100;
	13'd7720: q = 3'b100;
	13'd7721: q = 3'b100;
	13'd7722: q = 3'b100;
	13'd7723: q = 3'b100;
	13'd7724: q = 3'b100;
	13'd7725: q = 3'b100;
	13'd7726: q = 3'b100;
	13'd7727: q = 3'b100;
	13'd7728: q = 3'b100;
	13'd7729: q = 3'b100;
	13'd7730: q = 3'b100;
	13'd7731: q = 3'b100;
	13'd7732: q = 3'b100;
	13'd7733: q = 3'b100;
	13'd7734: q = 3'b100;
	13'd7735: q = 3'b100;
	13'd7736: q = 3'b100;
	13'd7737: q = 3'b100;
	13'd7738: q = 3'b100;
	13'd7739: q = 3'b100;
	13'd7740: q = 3'b100;
	13'd7741: q = 3'b100;
	13'd7742: q = 3'b100;
	13'd7743: q = 3'b100;
	13'd7744: q = 3'b100;
	13'd7745: q = 3'b100;
	13'd7746: q = 3'b100;
	13'd7747: q = 3'b100;
	13'd7748: q = 3'b100;
	13'd7749: q = 3'b100;
	13'd7750: q = 3'b100;
	13'd7751: q = 3'b100;
	13'd7752: q = 3'b100;
	13'd7753: q = 3'b100;
	13'd7754: q = 3'b100;
	13'd7755: q = 3'b100;
	13'd7756: q = 3'b100;
	13'd7757: q = 3'b100;
	13'd7758: q = 3'b100;
	13'd7759: q = 3'b100;
	13'd7760: q = 3'b100;
	13'd7761: q = 3'b100;
	13'd7762: q = 3'b100;
	13'd7763: q = 3'b100;
	13'd7764: q = 3'b100;
	13'd7765: q = 3'b100;
	13'd7766: q = 3'b100;
	13'd7767: q = 3'b100;
	13'd7768: q = 3'b100;
	13'd7769: q = 3'b100;
	13'd7770: q = 3'b100;
	13'd7771: q = 3'b100;
	13'd7772: q = 3'b100;
	13'd7773: q = 3'b100;
	13'd7774: q = 3'b100;
	13'd7775: q = 3'b100;
	13'd7776: q = 3'b100;
	13'd7777: q = 3'b100;
	13'd7778: q = 3'b100;
	13'd7779: q = 3'b100;
	13'd7780: q = 3'b100;
	13'd7781: q = 3'b100;
	13'd7782: q = 3'b100;
	13'd7783: q = 3'b100;
	13'd7784: q = 3'b100;
	13'd7785: q = 3'b100;
	13'd7786: q = 3'b100;
	13'd7787: q = 3'b100;
	13'd7788: q = 3'b100;
	13'd7789: q = 3'b100;
	13'd7790: q = 3'b100;
	13'd7791: q = 3'b100;
	13'd7792: q = 3'b100;
	13'd7793: q = 3'b100;
	13'd7794: q = 3'b100;
	13'd7795: q = 3'b100;
	13'd7796: q = 3'b100;
	13'd7797: q = 3'b100;
	13'd7798: q = 3'b100;
	13'd7799: q = 3'b100;
	13'd7800: q = 3'b100;
	13'd7801: q = 3'b100;
	13'd7802: q = 3'b100;
	13'd7803: q = 3'b100;
	13'd7804: q = 3'b100;
	13'd7805: q = 3'b100;
	13'd7806: q = 3'b100;
	13'd7807: q = 3'b100;
	13'd7808: q = 3'b100;
	13'd7809: q = 3'b100;
	13'd7810: q = 3'b100;
	13'd7811: q = 3'b100;
	13'd7812: q = 3'b100;
	13'd7813: q = 3'b100;
	13'd7814: q = 3'b100;
	13'd7815: q = 3'b100;
	13'd7816: q = 3'b100;
	13'd7817: q = 3'b100;
	13'd7818: q = 3'b100;
	13'd7819: q = 3'b100;
	13'd7820: q = 3'b100;
	13'd7821: q = 3'b100;
	13'd7822: q = 3'b100;
	13'd7823: q = 3'b100;
	13'd7824: q = 3'b100;
	13'd7825: q = 3'b100;
	13'd7826: q = 3'b100;
	13'd7827: q = 3'b100;
	13'd7828: q = 3'b100;
	13'd7829: q = 3'b100;
	13'd7830: q = 3'b100;
	13'd7831: q = 3'b100;
	13'd7832: q = 3'b100;
	13'd7833: q = 3'b100;
	13'd7834: q = 3'b100;
	13'd7835: q = 3'b100;
	13'd7836: q = 3'b100;
	13'd7837: q = 3'b100;
	13'd7838: q = 3'b100;
	13'd7839: q = 3'b100;
	13'd7840: q = 3'b100;
	13'd7841: q = 3'b100;
	13'd7842: q = 3'b100;
	13'd7843: q = 3'b100;
	13'd7844: q = 3'b100;
	13'd7845: q = 3'b100;
	13'd7846: q = 3'b100;
	13'd7847: q = 3'b100;
	13'd7848: q = 3'b100;
	13'd7849: q = 3'b100;
	13'd7850: q = 3'b100;
	13'd7851: q = 3'b100;
	13'd7852: q = 3'b100;
	13'd7853: q = 3'b100;
	13'd7854: q = 3'b100;
	13'd7855: q = 3'b100;
	13'd7856: q = 3'b100;
	13'd7857: q = 3'b100;
	13'd7858: q = 3'b100;
	13'd7859: q = 3'b100;
	13'd7860: q = 3'b100;
	13'd7861: q = 3'b100;
	13'd7862: q = 3'b100;
	13'd7863: q = 3'b100;
	13'd7864: q = 3'b100;
	13'd7865: q = 3'b100;
	13'd7866: q = 3'b100;
	13'd7867: q = 3'b100;
	13'd7868: q = 3'b100;
	13'd7869: q = 3'b100;
	13'd7870: q = 3'b100;
	13'd7871: q = 3'b100;
	13'd7872: q = 3'b000;
	13'd7873: q = 3'b000;
	13'd7874: q = 3'b100;
	13'd7875: q = 3'b100;
	13'd7876: q = 3'b100;
	13'd7877: q = 3'b100;
	13'd7878: q = 3'b100;
	13'd7879: q = 3'b100;
	13'd7880: q = 3'b100;
	13'd7881: q = 3'b100;
	13'd7882: q = 3'b100;
	13'd7883: q = 3'b100;
	13'd7884: q = 3'b100;
	13'd7885: q = 3'b100;
	13'd7886: q = 3'b100;
	13'd7887: q = 3'b100;
	13'd7888: q = 3'b100;
	13'd7889: q = 3'b100;
	13'd7890: q = 3'b100;
	13'd7891: q = 3'b100;
	13'd7892: q = 3'b100;
	13'd7893: q = 3'b100;
	13'd7894: q = 3'b100;
	13'd7895: q = 3'b100;
	13'd7896: q = 3'b100;
	13'd7897: q = 3'b100;
	13'd7898: q = 3'b100;
	13'd7899: q = 3'b100;
	13'd7900: q = 3'b100;
	13'd7901: q = 3'b100;
	13'd7902: q = 3'b000;
	13'd7903: q = 3'b000;
	13'd7904: q = 3'b000;
	13'd7905: q = 3'b000;
	13'd7906: q = 3'b100;
	13'd7907: q = 3'b100;
	13'd7908: q = 3'b100;
	13'd7909: q = 3'b100;
	13'd7910: q = 3'b100;
	13'd7911: q = 3'b100;
	13'd7912: q = 3'b100;
	13'd7913: q = 3'b100;
	13'd7914: q = 3'b100;
	13'd7915: q = 3'b100;
	13'd7916: q = 3'b100;
	13'd7917: q = 3'b100;
	13'd7918: q = 3'b100;
	13'd7919: q = 3'b100;
	13'd7920: q = 3'b100;
	13'd7921: q = 3'b100;
	13'd7922: q = 3'b100;
	13'd7923: q = 3'b100;
	13'd7924: q = 3'b100;
	13'd7925: q = 3'b100;
	13'd7926: q = 3'b100;
	13'd7927: q = 3'b100;
	13'd7928: q = 3'b100;
	13'd7929: q = 3'b100;
	13'd7930: q = 3'b100;
	13'd7931: q = 3'b100;
	13'd7932: q = 3'b100;
	13'd7933: q = 3'b100;
	13'd7934: q = 3'b000;
	13'd7935: q = 3'b000;
	13'd7936: q = 3'b000;
	13'd7937: q = 3'b000;
	13'd7938: q = 3'b100;
	13'd7939: q = 3'b100;
	13'd7940: q = 3'b100;
	13'd7941: q = 3'b100;
	13'd7942: q = 3'b100;
	13'd7943: q = 3'b100;
	13'd7944: q = 3'b100;
	13'd7945: q = 3'b100;
	13'd7946: q = 3'b100;
	13'd7947: q = 3'b100;
	13'd7948: q = 3'b100;
	13'd7949: q = 3'b100;
	13'd7950: q = 3'b100;
	13'd7951: q = 3'b100;
	13'd7952: q = 3'b100;
	13'd7953: q = 3'b100;
	13'd7954: q = 3'b100;
	13'd7955: q = 3'b100;
	13'd7956: q = 3'b100;
	13'd7957: q = 3'b100;
	13'd7958: q = 3'b100;
	13'd7959: q = 3'b100;
	13'd7960: q = 3'b100;
	13'd7961: q = 3'b100;
	13'd7962: q = 3'b100;
	13'd7963: q = 3'b100;
	13'd7964: q = 3'b100;
	13'd7965: q = 3'b100;
	13'd7966: q = 3'b000;
	13'd7967: q = 3'b000;
	13'd7968: q = 3'b000;
	13'd7969: q = 3'b000;
	13'd7970: q = 3'b100;
	13'd7971: q = 3'b100;
	13'd7972: q = 3'b100;
	13'd7973: q = 3'b100;
	13'd7974: q = 3'b100;
	13'd7975: q = 3'b100;
	13'd7976: q = 3'b100;
	13'd7977: q = 3'b100;
	13'd7978: q = 3'b100;
	13'd7979: q = 3'b100;
	13'd7980: q = 3'b100;
	13'd7981: q = 3'b100;
	13'd7982: q = 3'b100;
	13'd7983: q = 3'b100;
	13'd7984: q = 3'b100;
	13'd7985: q = 3'b100;
	13'd7986: q = 3'b100;
	13'd7987: q = 3'b100;
	13'd7988: q = 3'b100;
	13'd7989: q = 3'b100;
	13'd7990: q = 3'b100;
	13'd7991: q = 3'b100;
	13'd7992: q = 3'b100;
	13'd7993: q = 3'b100;
	13'd7994: q = 3'b100;
	13'd7995: q = 3'b100;
	13'd7996: q = 3'b100;
	13'd7997: q = 3'b100;
	13'd7998: q = 3'b000;
	13'd7999: q = 3'b000;
	13'd8000: q = 3'b000;
	13'd8001: q = 3'b000;
	13'd8002: q = 3'b000;
	13'd8003: q = 3'b000;
	13'd8004: q = 3'b100;
	13'd8005: q = 3'b100;
	13'd8006: q = 3'b100;
	13'd8007: q = 3'b100;
	13'd8008: q = 3'b100;
	13'd8009: q = 3'b100;
	13'd8010: q = 3'b100;
	13'd8011: q = 3'b100;
	13'd8012: q = 3'b100;
	13'd8013: q = 3'b100;
	13'd8014: q = 3'b100;
	13'd8015: q = 3'b100;
	13'd8016: q = 3'b100;
	13'd8017: q = 3'b100;
	13'd8018: q = 3'b100;
	13'd8019: q = 3'b100;
	13'd8020: q = 3'b100;
	13'd8021: q = 3'b100;
	13'd8022: q = 3'b100;
	13'd8023: q = 3'b100;
	13'd8024: q = 3'b100;
	13'd8025: q = 3'b100;
	13'd8026: q = 3'b100;
	13'd8027: q = 3'b100;
	13'd8028: q = 3'b000;
	13'd8029: q = 3'b000;
	13'd8030: q = 3'b000;
	13'd8031: q = 3'b000;
	13'd8032: q = 3'b000;
	13'd8033: q = 3'b000;
	13'd8034: q = 3'b000;
	13'd8035: q = 3'b000;
	13'd8036: q = 3'b100;
	13'd8037: q = 3'b100;
	13'd8038: q = 3'b100;
	13'd8039: q = 3'b100;
	13'd8040: q = 3'b100;
	13'd8041: q = 3'b100;
	13'd8042: q = 3'b100;
	13'd8043: q = 3'b100;
	13'd8044: q = 3'b100;
	13'd8045: q = 3'b100;
	13'd8046: q = 3'b100;
	13'd8047: q = 3'b100;
	13'd8048: q = 3'b100;
	13'd8049: q = 3'b100;
	13'd8050: q = 3'b100;
	13'd8051: q = 3'b100;
	13'd8052: q = 3'b100;
	13'd8053: q = 3'b100;
	13'd8054: q = 3'b100;
	13'd8055: q = 3'b100;
	13'd8056: q = 3'b100;
	13'd8057: q = 3'b100;
	13'd8058: q = 3'b100;
	13'd8059: q = 3'b100;
	13'd8060: q = 3'b000;
	13'd8061: q = 3'b000;
	13'd8062: q = 3'b000;
	13'd8063: q = 3'b000;
	13'd8064: q = 3'b000;
	13'd8065: q = 3'b000;
	13'd8066: q = 3'b000;
	13'd8067: q = 3'b000;
	13'd8068: q = 3'b000;
	13'd8069: q = 3'b000;
	13'd8070: q = 3'b100;
	13'd8071: q = 3'b100;
	13'd8072: q = 3'b100;
	13'd8073: q = 3'b100;
	13'd8074: q = 3'b100;
	13'd8075: q = 3'b100;
	13'd8076: q = 3'b100;
	13'd8077: q = 3'b100;
	13'd8078: q = 3'b100;
	13'd8079: q = 3'b100;
	13'd8080: q = 3'b100;
	13'd8081: q = 3'b100;
	13'd8082: q = 3'b100;
	13'd8083: q = 3'b100;
	13'd8084: q = 3'b100;
	13'd8085: q = 3'b100;
	13'd8086: q = 3'b100;
	13'd8087: q = 3'b100;
	13'd8088: q = 3'b100;
	13'd8089: q = 3'b100;
	13'd8090: q = 3'b000;
	13'd8091: q = 3'b000;
	13'd8092: q = 3'b000;
	13'd8093: q = 3'b000;
	13'd8094: q = 3'b000;
	13'd8095: q = 3'b000;
	13'd8096: q = 3'b000;
	13'd8097: q = 3'b000;
	13'd8098: q = 3'b000;
	13'd8099: q = 3'b000;
	13'd8100: q = 3'b000;
	13'd8101: q = 3'b000;
	13'd8102: q = 3'b100;
	13'd8103: q = 3'b100;
	13'd8104: q = 3'b100;
	13'd8105: q = 3'b100;
	13'd8106: q = 3'b100;
	13'd8107: q = 3'b100;
	13'd8108: q = 3'b100;
	13'd8109: q = 3'b100;
	13'd8110: q = 3'b100;
	13'd8111: q = 3'b100;
	13'd8112: q = 3'b100;
	13'd8113: q = 3'b100;
	13'd8114: q = 3'b100;
	13'd8115: q = 3'b100;
	13'd8116: q = 3'b100;
	13'd8117: q = 3'b100;
	13'd8118: q = 3'b100;
	13'd8119: q = 3'b100;
	13'd8120: q = 3'b100;
	13'd8121: q = 3'b100;
	13'd8122: q = 3'b000;
	13'd8123: q = 3'b000;
	13'd8124: q = 3'b000;
	13'd8125: q = 3'b000;
	13'd8126: q = 3'b000;
	13'd8127: q = 3'b000;
	13'd8128: q = 3'b000;
	13'd8129: q = 3'b000;
	13'd8130: q = 3'b000;
	13'd8131: q = 3'b000;
	13'd8132: q = 3'b000;
	13'd8133: q = 3'b000;
	13'd8134: q = 3'b000;
	13'd8135: q = 3'b000;
	13'd8136: q = 3'b000;
	13'd8137: q = 3'b000;
	13'd8138: q = 3'b100;
	13'd8139: q = 3'b100;
	13'd8140: q = 3'b100;
	13'd8141: q = 3'b100;
	13'd8142: q = 3'b100;
	13'd8143: q = 3'b100;
	13'd8144: q = 3'b100;
	13'd8145: q = 3'b100;
	13'd8146: q = 3'b100;
	13'd8147: q = 3'b100;
	13'd8148: q = 3'b100;
	13'd8149: q = 3'b100;
	13'd8150: q = 3'b000;
	13'd8151: q = 3'b000;
	13'd8152: q = 3'b000;
	13'd8153: q = 3'b000;
	13'd8154: q = 3'b000;
	13'd8155: q = 3'b000;
	13'd8156: q = 3'b000;
	13'd8157: q = 3'b000;
	13'd8158: q = 3'b000;
	13'd8159: q = 3'b000;
	13'd8160: q = 3'b000;
	13'd8161: q = 3'b000;
	13'd8162: q = 3'b000;
	13'd8163: q = 3'b000;
	13'd8164: q = 3'b000;
	13'd8165: q = 3'b000;
	13'd8166: q = 3'b000;
	13'd8167: q = 3'b000;
	13'd8168: q = 3'b000;
	13'd8169: q = 3'b000;
	13'd8170: q = 3'b100;
	13'd8171: q = 3'b100;
	13'd8172: q = 3'b100;
	13'd8173: q = 3'b100;
	13'd8174: q = 3'b100;
	13'd8175: q = 3'b100;
	13'd8176: q = 3'b100;
	13'd8177: q = 3'b100;
	13'd8178: q = 3'b100;
	13'd8179: q = 3'b100;
	13'd8180: q = 3'b100;
	13'd8181: q = 3'b100;
	13'd8182: q = 3'b000;
	13'd8183: q = 3'b000;
	13'd8184: q = 3'b000;
	13'd8185: q = 3'b000;
	13'd8186: q = 3'b000;
	13'd8187: q = 3'b000;
	13'd8188: q = 3'b000;
	13'd8189: q = 3'b000;
	13'd8190: q = 3'b000;
	13'd8191: q = 3'b000;
	endcase

endmodule

